CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1278 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 450 89 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3675 0 0
2
43488.4 0
0
13 Logic Switch~
5 325 88 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7278 0 0
2
43488.4 0
0
13 Logic Switch~
5 201 89 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
926 0 0
2
43488.4 0
0
13 Logic Switch~
5 75 86 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -22 9 -14
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6747 0 0
2
43488.4 0
0
7 Ground~
168 1183 44 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5177 0 0
2
43488.4 0
0
9 CC 7-Seg~
183 1186 123 0 17 19
10 9 8 7 6 5 4 3 35 2
1 1 1 1 0 1 1 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
5594 0 0
2
43488.4 0
0
8 2-In OR~
219 786 887 0 3 22
0 11 10 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
9933 0 0
2
43488.4 0
0
8 2-In OR~
219 687 840 0 3 22
0 13 12 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
8987 0 0
2
43488.4 0
0
6 74136~
219 580 873 0 3 22
0 15 14 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U10A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3275 0 0
2
43488.4 0
0
9 2-In AND~
219 591 820 0 3 22
0 14 16 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3551 0 0
2
43488.4 0
0
8 2-In OR~
219 781 723 0 3 22
0 18 17 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
9522 0 0
2
43488.4 0
0
9 2-In AND~
219 697 769 0 3 22
0 19 15 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3443 0 0
2
43488.4 0
0
8 2-In OR~
219 586 756 0 3 22
0 20 16 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3935 0 0
2
43488.4 0
0
8 2-In OR~
219 700 666 0 3 22
0 10 21 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
4532 0 0
2
43488.4 0
0
9 2-In AND~
219 593 700 0 3 22
0 20 16 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7600 0 0
2
43488.4 0
0
9 2-In AND~
219 696 587 0 3 22
0 22 16 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
6952 0 0
2
43488.4 0
0
8 2-In OR~
219 583 577 0 3 22
0 23 14 22
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3663 0 0
2
43488.4 0
0
8 2-In OR~
219 920 503 0 3 22
0 25 24 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9511 0 0
2
43488.4 0
0
5 7415~
219 595 520 0 4 22
0 15 20 26 24
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
4625 0 0
2
43488.4 0
0
9 2-In AND~
219 596 477 0 3 22
0 14 16 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
6215 0 0
2
43488.4 0
0
8 2-In OR~
219 831 463 0 3 22
0 28 27 25
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4535 0 0
2
43488.4 0
0
9 2-In AND~
219 761 437 0 3 22
0 29 23 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3611 0 0
2
43488.4 0
0
8 2-In OR~
219 679 423 0 3 22
0 30 16 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9183 0 0
2
43488.4 0
0
8 2-In OR~
219 592 408 0 3 22
0 10 14 30
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3593 0 0
2
43488.4 0
0
8 2-In OR~
219 669 348 0 3 22
0 31 26 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4142 0 0
2
43488.4 0
0
8 2-In OR~
219 594 337 0 3 22
0 15 20 31
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9564 0 0
2
43488.4 0
0
8 2-In OR~
219 670 279 0 3 22
0 32 23 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7772 0 0
2
43488.4 0
0
6 74266~
219 594 268 0 3 22
0 14 26 32
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3826 0 0
2
43488.4 0
0
8 2-In OR~
219 746 204 0 3 22
0 33 10 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9216 0 0
2
43488.4 0
0
8 2-In OR~
219 666 195 0 3 22
0 34 14 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
770 0 0
2
43488.4 0
0
6 74266~
219 588 187 0 3 22
0 15 26 34
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6894 0 0
2
43488.4 0
0
9 Inverter~
13 497 140 0 2 22
0 26 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3840 0 0
2
43488.4 0
0
9 Inverter~
13 372 142 0 2 22
0 14 20
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
6568 0 0
2
43488.4 0
0
9 Inverter~
13 247 143 0 2 22
0 15 23
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
656 0 0
2
43488.4 0
0
62
1 9 2 0 0 8320 0 5 6 0 0 3
1183 52
1186 52
1186 81
3 7 3 0 0 8320 0 7 6 0 0 3
819 887
1201 887
1201 159
3 6 4 0 0 8320 0 11 6 0 0 3
814 723
1195 723
1195 159
3 5 5 0 0 4224 0 16 6 0 0 3
717 587
1189 587
1189 159
3 4 6 0 0 8320 0 18 6 0 0 3
953 503
1183 503
1183 159
3 3 7 0 0 4224 0 25 6 0 0 3
702 348
1177 348
1177 159
3 2 8 0 0 4224 0 27 6 0 0 3
703 279
1171 279
1171 159
3 1 9 0 0 4224 0 29 6 0 0 3
779 204
1165 204
1165 159
0 2 10 0 0 8320 0 0 7 24 0 3
75 656
75 896
773 896
3 1 11 0 0 8320 0 8 7 0 0 3
720 840
720 878
773 878
3 2 12 0 0 4224 0 9 8 0 0 3
613 873
674 873
674 849
3 1 13 0 0 4224 0 10 8 0 0 3
612 820
674 820
674 831
0 2 14 0 0 8192 0 0 9 16 0 3
325 811
325 882
564 882
0 1 15 0 0 8192 0 0 9 19 0 3
201 777
201 864
564 864
0 2 16 0 0 8192 0 0 10 21 0 3
500 765
500 829
567 829
0 1 14 0 0 8192 0 0 10 29 0 3
325 584
325 811
567 811
3 2 17 0 0 4224 0 12 11 0 0 3
718 769
768 769
768 732
3 1 18 0 0 4224 0 14 11 0 0 3
733 666
733 714
768 714
0 2 15 0 0 8320 0 0 12 35 0 3
201 511
201 778
673 778
3 1 19 0 0 4224 0 13 12 0 0 3
619 756
673 756
673 760
0 2 16 0 0 8192 0 0 13 25 0 3
500 709
500 765
573 765
0 1 20 0 0 8192 0 0 13 26 0 3
375 691
375 747
573 747
3 2 21 0 0 4224 0 15 14 0 0 3
614 700
687 700
687 675
0 1 10 0 0 0 0 0 14 45 0 3
75 399
75 657
687 657
0 2 16 0 0 4096 0 0 15 27 0 3
500 596
500 709
569 709
0 1 20 0 0 0 0 0 15 34 0 3
375 520
375 691
569 691
0 2 16 0 0 8192 0 0 16 38 0 3
500 483
500 596
672 596
3 1 22 0 0 8320 0 17 16 0 0 3
616 577
616 578
672 578
0 2 14 0 0 8192 0 0 17 39 0 3
325 468
325 586
570 586
0 1 23 0 0 8192 0 0 17 40 0 3
250 446
250 568
570 568
4 2 24 0 0 4224 0 19 18 0 0 3
616 520
907 520
907 512
3 1 25 0 0 4224 0 21 18 0 0 3
864 463
907 463
907 494
0 3 26 0 0 4096 0 0 19 46 0 3
450 357
450 529
571 529
0 2 20 0 0 0 0 0 19 48 0 3
375 345
375 520
571 520
0 1 15 0 0 0 0 0 19 49 0 3
201 328
201 511
571 511
3 2 27 0 0 4224 0 20 21 0 0 3
617 477
818 477
818 472
3 1 28 0 0 4224 0 22 21 0 0 3
782 437
818 437
818 454
0 2 16 0 0 0 0 0 20 42 0 3
500 431
500 486
572 486
0 1 14 0 0 8192 0 0 20 44 0 3
325 417
325 468
572 468
0 2 23 0 0 8320 0 0 22 50 0 3
250 288
250 446
737 446
3 1 29 0 0 4224 0 23 22 0 0 3
712 423
737 423
737 428
2 2 16 0 0 4224 0 32 23 0 0 3
500 158
500 432
666 432
3 1 30 0 0 4224 0 24 23 0 0 3
625 408
666 408
666 414
0 2 14 0 0 8192 0 0 24 53 0 3
325 259
325 417
579 417
0 1 10 0 0 0 0 0 24 54 0 3
75 212
75 399
579 399
0 2 26 0 0 8320 0 0 25 52 0 3
450 277
450 357
656 357
3 1 31 0 0 8320 0 26 25 0 0 3
627 337
627 339
656 339
2 2 20 0 0 8320 0 33 26 0 0 3
375 160
375 346
581 346
0 1 15 0 0 0 0 0 26 59 0 3
201 177
201 328
581 328
2 2 23 0 0 0 0 34 27 0 0 3
250 161
250 288
657 288
3 1 32 0 0 4224 0 28 27 0 0 4
633 268
645 268
645 270
657 270
0 2 26 0 0 0 0 0 28 58 0 3
450 195
450 277
578 277
0 1 14 0 0 0 0 0 28 56 0 3
325 203
325 259
578 259
1 2 10 0 0 0 0 4 29 0 0 3
75 98
75 213
733 213
3 1 33 0 0 4224 0 30 29 0 0 2
699 195
733 195
1 2 14 0 0 8320 0 2 30 0 0 3
325 100
325 204
653 204
3 1 34 0 0 8320 0 31 30 0 0 3
627 187
627 186
653 186
1 2 26 0 0 0 0 1 31 0 0 3
450 101
450 196
572 196
1 1 15 0 0 0 0 3 31 0 0 3
201 101
201 178
572 178
1 1 26 0 0 0 0 1 32 0 0 3
450 101
500 101
500 122
1 1 14 0 0 0 0 2 33 0 0 3
325 100
375 100
375 124
1 1 15 0 0 0 0 3 34 0 0 3
201 101
250 101
250 125
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
431 11 469 26
446 23 453 34
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
306 12 342 27
320 24 327 35
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
183 13 219 28
197 24 204 35
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
57 11 95 26
72 23 79 34
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
