CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
76546066 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 406 52 0 1 11
0 25
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9265 0 0
2
43490.3 0
0
13 Logic Switch~
5 298 51 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
43490.3 1
0
13 Logic Switch~
5 175 63 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
43490.3 2
0
13 Logic Switch~
5 45 68 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9968 0 0
2
43490.3 3
0
14 Logic Display~
6 963 359 0 1 2
10 34
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
9281 0 0
2
5.89878e-315 0
0
7 Ground~
168 1098 153 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8464 0 0
2
5.89878e-315 0
0
9 CC 7-Seg~
183 848 75 0 17 19
10 9 8 7 6 5 4 3 35 2
1 1 1 0 0 1 1 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7168 0 0
2
43490.3 4
0
8 2-In OR~
219 661 568 0 3 22
0 11 10 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3171 0 0
2
43490.3 5
0
6 74136~
219 524 592 0 3 22
0 14 13 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4139 0 0
2
43490.3 6
0
8 2-In OR~
219 585 549 0 3 22
0 15 12 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
6435 0 0
2
43490.3 7
0
9 2-In AND~
219 516 545 0 3 22
0 13 16 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
5283 0 0
2
43490.3 8
0
8 2-In OR~
219 666 475 0 3 22
0 18 17 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
6874 0 0
2
43490.3 9
0
9 2-In AND~
219 594 499 0 3 22
0 19 14 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
5305 0 0
2
43490.3 10
0
8 2-In OR~
219 510 491 0 3 22
0 20 16 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
34 0 0
2
43490.3 11
0
8 2-In OR~
219 576 451 0 3 22
0 21 10 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
969 0 0
2
43490.3 12
0
9 2-In AND~
219 520 444 0 3 22
0 20 16 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
8402 0 0
2
43490.3 13
0
9 2-In AND~
219 594 403 0 3 22
0 22 16 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3751 0 0
2
43490.3 14
0
8 2-In OR~
219 513 391 0 3 22
0 23 13 22
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4292 0 0
2
43490.3 15
0
5 7415~
219 523 349 0 4 22
0 14 20 25 24
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 7 0
1 U
6118 0 0
2
43490.3 16
0
9 2-In AND~
219 516 314 0 3 22
0 13 16 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
34 0 0
2
43490.3 17
0
8 3-In OR~
219 648 270 0 4 22
0 27 26 24 6
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
6357 0 0
2
43490.3 18
0
9 2-In AND~
219 592 241 0 3 22
0 28 23 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
319 0 0
2
43490.3 19
0
8 3-In OR~
219 504 244 0 4 22
0 10 13 16 28
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 3 0
1 U
3976 0 0
2
43490.3 20
0
8 3-In OR~
219 503 199 0 4 22
0 14 20 25 7
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 3 0
1 U
7634 0 0
2
43490.3 21
0
8 2-In OR~
219 634 134 0 3 22
0 29 23 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
523 0 0
2
43490.3 22
0
9 Inverter~
13 586 112 0 2 22
0 30 29
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
6748 0 0
2
43490.3 23
0
6 74136~
219 531 126 0 3 22
0 13 25 30
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6901 0 0
2
43490.3 24
0
8 3-In OR~
219 697 52 0 4 22
0 31 10 13 9
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
842 0 0
2
43490.3 25
0
9 Inverter~
13 584 77 0 2 22
0 32 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3277 0 0
2
43490.3 26
0
6 74136~
219 532 75 0 3 22
0 14 25 32
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4212 0 0
2
43490.3 27
0
9 Inverter~
13 437 110 0 2 22
0 25 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
4720 0 0
2
43490.3 36
0
9 Inverter~
13 337 114 0 2 22
0 13 20
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
5551 0 0
2
43490.3 37
0
9 Inverter~
13 231 114 0 2 22
0 14 23
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
6986 0 0
2
43490.3 38
0
9 Inverter~
13 91 107 0 2 22
0 10 33
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8745 0 0
2
43490.3 39
0
69
9 1 2 0 0 8320 0 7 6 0 0 4
848 33
848 29
1098 29
1098 147
7 3 3 0 0 4224 0 7 8 0 0 3
863 111
863 568
694 568
3 6 4 0 0 8320 0 12 7 0 0 3
699 475
857 475
857 111
5 3 5 0 0 4224 0 7 17 0 0 3
851 111
851 403
615 403
4 4 6 0 0 16512 0 21 7 0 0 5
681 270
734 270
734 276
845 276
845 111
4 3 7 0 0 12416 0 24 7 0 0 5
536 199
684 199
684 206
839 206
839 111
3 2 8 0 0 12416 0 25 7 0 0 7
667 134
683 134
683 135
792 135
792 175
833 175
833 111
4 1 9 0 0 8320 0 28 7 0 0 5
730 52
796 52
796 170
827 170
827 111
0 2 10 0 0 4224 0 0 8 69 0 4
45 572
627 572
627 577
648 577
3 1 11 0 0 4224 0 10 8 0 0 4
618 549
633 549
633 559
648 559
3 2 12 0 0 8320 0 9 10 0 0 4
557 592
555 592
555 558
572 558
0 2 13 0 0 4096 0 0 9 65 0 4
298 575
494 575
494 601
508 601
0 1 14 0 0 4096 0 0 9 67 0 2
175 583
508 583
3 1 15 0 0 12416 0 11 10 0 0 4
537 545
553 545
553 540
572 540
0 2 16 0 0 4096 0 0 11 62 0 2
439 554
492 554
0 1 13 0 0 0 0 0 11 65 0 2
298 536
492 536
3 2 17 0 0 4224 0 13 12 0 0 4
615 499
635 499
635 484
653 484
3 1 18 0 0 4224 0 15 12 0 0 4
609 451
635 451
635 466
653 466
0 2 14 0 0 4096 0 0 13 67 0 4
175 515
552 515
552 508
570 508
3 1 19 0 0 12416 0 14 13 0 0 4
543 491
552 491
552 490
570 490
0 2 16 0 0 0 0 0 14 62 0 4
439 504
454 504
454 500
497 500
0 1 20 0 0 12288 0 0 14 64 0 4
340 486
355 486
355 482
497 482
0 2 10 0 0 0 0 0 15 69 0 4
45 465
551 465
551 460
563 460
3 1 21 0 0 12416 0 16 15 0 0 4
541 444
551 444
551 442
563 442
0 2 16 0 0 0 0 0 16 62 0 4
439 454
454 454
454 453
496 453
0 1 20 0 0 0 0 0 16 64 0 4
340 436
355 436
355 435
496 435
0 2 16 0 0 4096 0 0 17 62 0 4
439 420
556 420
556 412
570 412
3 1 22 0 0 12416 0 18 17 0 0 4
546 391
556 391
556 394
570 394
0 2 13 0 0 0 0 0 18 65 0 4
298 404
492 404
492 400
500 400
0 1 23 0 0 12288 0 0 18 66 0 4
234 385
249 385
249 382
500 382
4 3 24 0 0 4224 0 19 21 0 0 4
544 349
620 349
620 279
635 279
0 3 25 0 0 4096 0 0 19 63 0 4
406 362
487 362
487 358
499 358
0 2 20 0 0 12288 0 0 19 64 0 4
340 352
355 352
355 349
499 349
0 1 14 0 0 0 0 0 19 67 0 4
175 343
190 343
190 340
499 340
3 2 26 0 0 4224 0 20 21 0 0 4
537 314
625 314
625 270
636 270
0 2 16 0 0 0 0 0 20 62 0 2
439 323
492 323
0 1 13 0 0 0 0 0 20 65 0 2
298 305
492 305
3 1 27 0 0 8320 0 22 21 0 0 4
613 241
625 241
625 261
635 261
0 2 23 0 0 4096 0 0 22 66 0 4
234 283
561 283
561 250
568 250
4 1 28 0 0 4224 0 23 22 0 0 4
537 244
561 244
561 232
568 232
0 3 16 0 0 0 0 0 23 62 0 4
439 269
454 269
454 253
491 253
0 2 13 0 0 0 0 0 23 65 0 4
298 260
313 260
313 244
492 244
0 1 10 0 0 0 0 0 23 69 0 4
45 251
60 251
60 235
491 235
0 3 25 0 0 0 0 0 24 63 0 4
406 215
421 215
421 208
490 208
0 2 20 0 0 0 0 0 24 64 0 4
340 206
355 206
355 199
491 199
0 1 14 0 0 0 0 0 24 67 0 4
175 197
190 197
190 190
490 190
0 2 23 0 0 4096 0 0 25 66 0 4
234 168
611 168
611 143
621 143
2 1 29 0 0 8320 0 26 25 0 0 4
607 112
611 112
611 125
621 125
3 1 30 0 0 8320 0 27 26 0 0 4
564 126
558 126
558 112
571 112
0 2 25 0 0 12288 0 0 27 63 0 4
406 140
421 140
421 135
515 135
0 1 13 0 0 0 0 0 27 65 0 4
298 139
493 139
493 117
515 117
0 3 13 0 0 0 0 0 28 65 0 6
298 81
494 81
494 47
610 47
610 61
684 61
0 2 10 0 0 0 0 0 28 69 0 6
45 121
77 121
77 35
610 35
610 52
685 52
2 1 31 0 0 12416 0 29 28 0 0 4
605 77
615 77
615 43
684 43
3 1 32 0 0 12416 0 30 29 0 0 4
565 75
562 75
562 77
569 77
0 2 25 0 0 0 0 0 30 58 0 3
438 82
438 84
516 84
0 1 14 0 0 0 0 0 30 60 0 5
212 91
212 68
490 68
490 66
516 66
0 1 25 0 0 0 0 0 31 63 0 3
406 82
440 82
440 92
0 1 13 0 0 0 0 0 32 65 0 3
298 83
340 83
340 96
0 1 14 0 0 0 0 0 33 67 0 3
175 91
234 91
234 96
0 1 10 0 0 0 0 0 34 69 0 3
45 90
94 90
94 89
2 0 16 0 0 12416 0 31 0 0 0 6
440 128
440 269
439 269
439 585
459 585
459 593
1 0 25 0 0 4224 0 1 0 0 0 4
406 64
406 586
393 586
393 594
2 0 20 0 0 4224 0 32 0 0 0 4
340 132
340 590
329 590
329 598
1 0 13 0 0 4224 0 2 0 0 0 4
298 63
298 593
273 593
273 601
2 0 23 0 0 4224 0 33 0 0 0 4
234 132
234 597
213 597
213 605
1 0 14 0 0 4224 0 3 0 0 0 4
175 75
175 594
148 594
148 602
2 0 33 0 0 4224 0 34 0 0 0 4
94 125
94 596
79 596
79 604
1 0 10 0 0 0 0 4 0 0 0 4
45 80
45 598
39 598
39 606
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
687 534 716 558
697 542 705 558
1 g
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
684 441 713 465
694 449 702 465
1 f
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
610 369 639 393
620 377 628 393
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
679 241 708 265
689 249 697 265
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
541 176 570 200
551 184 559 200
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
657 106 686 130
667 114 675 130
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
664 31 693 55
674 39 682 55
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
437 36 466 60
447 44 455 60
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
313 56 342 80
323 64 331 80
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
195 43 224 67
205 51 213 67
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
83 44 112 68
93 52 101 68
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
