CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
47
13 Logic Switch~
5 172 38 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 141 39 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 112 39 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 79 39 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 342 604 0 3 22
0 12 10 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
8157 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 262 595 0 3 22
0 14 13 12
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
5572 0 0
2
5.89878e-315 0
0
9 Inverter~
13 207 612 0 2 22
0 15 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
8901 0 0
2
5.89878e-315 0
0
9 Inverter~
13 204 581 0 2 22
0 16 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
7361 0 0
2
5.89878e-315 0
0
7 Ground~
168 884 158 0 1 3
0 2
0
0 0 53360 90
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
5.89878e-315 0
0
9 CC 7-Seg~
183 759 206 0 17 19
10 9 8 7 6 5 4 3 48 2
1 0 1 1 1 1 1 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 402 736 0 3 22
0 18 17 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3472 0 0
2
5.89878e-315 0
0
9 Inverter~
13 208 728 0 2 22
0 15 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
9998 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 264 719 0 3 22
0 16 19 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3536 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 317 680 0 3 22
0 21 20 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
4597 0 0
2
5.89878e-315 0
0
6 74136~
219 211 672 0 3 22
0 10 16 21
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3835 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 392 553 0 3 22
0 22 11 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3670 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 313 543 0 3 22
0 23 17 22
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
5616 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 264 523 0 3 22
0 25 24 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
9323 0 0
2
5.89878e-315 0
0
9 Inverter~
13 203 544 0 2 22
0 15 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 6 0
1 U
317 0 0
2
5.89878e-315 0
0
9 Inverter~
13 202 515 0 2 22
0 16 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
3108 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 402 466 0 3 22
0 27 26 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4299 0 0
2
5.89878e-315 0
0
9 Inverter~
13 204 482 0 2 22
0 15 26
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
9672 0 0
2
5.89878e-315 0
0
9 Inverter~
13 204 448 0 2 22
0 10 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
7876 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 248 457 0 3 22
0 28 16 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
6369 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 333 365 0 3 22
0 30 31 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9172 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 297 400 0 3 22
0 32 33 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7100 0 0
2
5.89878e-315 0
0
9 Inverter~
13 244 424 0 2 22
0 16 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
3820 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 210 393 0 3 22
0 10 15 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
7678 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 395 311 0 3 22
0 34 29 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
961 0 0
2
5.89878e-315 0
0
9 Inverter~
13 201 362 0 2 22
0 15 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
3178 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 273 353 0 3 22
0 16 35 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3409 0 0
2
5.89878e-315 0
0
9 Inverter~
13 201 319 0 2 22
0 10 36
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
3951 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 329 281 0 3 22
0 37 36 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8885 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 257 270 0 3 22
0 39 38 37
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3780 0 0
2
5.89878e-315 0
0
9 Inverter~
13 201 295 0 2 22
0 15 38
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
9265 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 199 262 0 3 22
0 17 16 39
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9442 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 396 212 0 3 22
0 40 15 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9424 0 0
2
5.89878e-315 0
0
9 Inverter~
13 197 214 0 2 22
0 16 41
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
9968 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 250 205 0 3 22
0 10 41 40
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9281 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 393 147 0 3 22
0 43 42 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8464 0 0
2
5.89878e-315 0
0
9 Inverter~
13 250 164 0 2 22
0 10 42
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
7168 0 0
2
5.89878e-315 0
0
9 Inverter~
13 250 137 0 2 22
0 44 43
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3171 0 0
2
5.89878e-315 0
0
6 74136~
219 200 138 0 3 22
0 16 15 44
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4139 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 308 100 0 3 22
0 46 17 45
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1B
-8 -27 13 -19
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6435 0 0
2
5.89878e-315 0
0
9 Inverter~
13 250 91 0 2 22
0 47 46
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
5283 0 0
2
5.89878e-315 0
0
6 74136~
219 198 91 0 3 22
0 10 15 47
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6874 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 393 63 0 3 22
0 16 45 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5305 0 0
2
5.89878e-315 0
0
80
1 9 2 0 0 4224 0 9 10 0 0 3
877 159
759 159
759 164
7 3 3 0 0 4224 0 10 11 0 0 3
774 242
774 736
435 736
6 3 4 0 0 8320 0 10 16 0 0 3
768 242
768 553
425 553
5 3 5 0 0 8320 0 10 21 0 0 3
762 242
762 466
423 466
4 3 6 0 0 8336 0 10 29 0 0 5
756 242
756 282
446 282
446 311
428 311
3 3 7 0 0 8320 0 10 37 0 0 5
750 242
750 270
472 270
472 212
429 212
2 3 8 0 0 8320 0 10 40 0 0 5
744 242
744 256
484 256
484 147
426 147
1 3 9 0 0 8320 0 10 47 0 0 5
738 242
738 246
495 246
495 63
426 63
0 2 10 0 0 4096 0 0 5 79 0 4
113 627
310 627
310 613
318 613
3 2 11 0 0 8320 0 5 16 0 0 4
363 604
371 604
371 562
379 562
3 1 12 0 0 4224 0 6 5 0 0 2
295 595
318 595
2 2 13 0 0 4224 0 7 6 0 0 4
228 612
241 612
241 604
249 604
2 1 14 0 0 4224 0 8 6 0 0 4
225 581
241 581
241 586
249 586
0 1 15 0 0 4096 0 0 7 77 0 2
172 612
192 612
0 1 16 0 0 4096 0 0 8 78 0 4
140 582
181 582
181 581
189 581
0 2 17 0 0 4096 0 0 11 80 0 2
78 745
389 745
3 1 18 0 0 8320 0 14 11 0 0 4
350 680
381 680
381 727
389 727
0 1 15 0 0 4096 0 0 12 77 0 2
172 728
193 728
2 2 19 0 0 4224 0 12 13 0 0 2
229 728
240 728
0 1 16 0 0 4096 0 0 13 78 0 2
140 710
240 710
3 2 20 0 0 8320 0 13 14 0 0 4
285 719
295 719
295 689
304 689
3 1 21 0 0 12416 0 15 14 0 0 4
244 672
251 672
251 671
304 671
0 2 16 0 0 0 0 0 15 78 0 4
140 682
187 682
187 681
195 681
0 1 10 0 0 0 0 0 15 79 0 2
113 663
195 663
3 1 22 0 0 12416 0 17 16 0 0 4
346 543
357 543
357 544
379 544
0 2 17 0 0 0 0 0 17 80 0 2
78 552
300 552
3 1 23 0 0 8320 0 18 17 0 0 4
285 523
292 523
292 534
300 534
2 2 24 0 0 8320 0 19 18 0 0 4
224 544
232 544
232 532
240 532
2 1 25 0 0 4224 0 20 18 0 0 4
223 515
232 515
232 514
240 514
0 1 15 0 0 0 0 0 19 77 0 2
172 544
188 544
0 1 16 0 0 0 0 0 20 78 0 4
140 516
179 516
179 515
187 515
2 2 26 0 0 4224 0 22 21 0 0 4
225 482
370 482
370 475
378 475
3 1 27 0 0 4224 0 24 21 0 0 2
281 457
378 457
0 1 15 0 0 0 0 0 22 77 0 2
171 482
189 482
0 1 10 0 0 0 0 0 23 79 0 2
113 448
189 448
2 1 28 0 0 4224 0 23 24 0 0 2
225 448
235 448
0 2 16 0 0 0 0 0 24 78 0 2
141 466
235 466
3 2 29 0 0 8320 0 25 29 0 0 6
366 365
370 365
370 330
361 330
361 320
382 320
3 1 30 0 0 4224 0 31 25 0 0 4
294 353
312 353
312 356
320 356
2 3 31 0 0 4224 0 25 26 0 0 3
320 374
320 400
318 400
3 1 32 0 0 4224 0 28 26 0 0 4
231 393
265 393
265 391
273 391
2 2 33 0 0 8320 0 27 26 0 0 4
265 424
269 424
269 409
273 409
0 1 16 0 0 0 0 0 27 78 0 2
141 424
229 424
0 2 15 0 0 0 0 0 28 77 0 4
172 403
178 403
178 402
186 402
0 1 10 0 0 0 0 0 28 79 0 2
113 384
186 384
3 1 34 0 0 12416 0 33 29 0 0 4
350 281
358 281
358 302
382 302
0 1 15 0 0 0 0 0 30 77 0 2
172 362
186 362
2 2 35 0 0 4224 0 30 31 0 0 2
222 362
249 362
0 1 16 0 0 4096 0 0 31 78 0 2
141 344
249 344
2 2 36 0 0 4224 0 32 33 0 0 4
222 319
297 319
297 290
305 290
0 1 10 0 0 0 0 0 32 79 0 2
113 319
186 319
3 1 37 0 0 12416 0 34 33 0 0 4
290 270
297 270
297 272
305 272
2 2 38 0 0 8320 0 35 34 0 0 4
222 295
236 295
236 279
244 279
3 1 39 0 0 12416 0 36 34 0 0 4
232 262
236 262
236 261
244 261
0 1 15 0 0 0 0 0 35 77 0 2
172 295
186 295
0 2 16 0 0 0 0 0 36 78 0 2
141 271
186 271
0 1 17 0 0 0 0 0 36 80 0 2
79 253
186 253
0 2 15 0 0 4096 0 0 37 77 0 4
172 229
375 229
375 221
383 221
3 1 40 0 0 4224 0 39 37 0 0 4
283 205
375 205
375 203
383 203
2 2 41 0 0 4224 0 38 39 0 0 2
218 214
237 214
0 1 16 0 0 0 0 0 38 78 0 2
141 214
182 214
0 1 10 0 0 0 0 0 39 79 0 2
113 196
237 196
0 2 15 0 0 0 0 0 43 77 0 2
172 147
184 147
2 2 42 0 0 4224 0 41 40 0 0 4
271 164
372 164
372 156
380 156
2 1 43 0 0 4224 0 42 40 0 0 4
271 137
372 137
372 138
380 138
0 1 10 0 0 0 0 0 41 79 0 2
113 164
235 164
3 1 44 0 0 8320 0 43 42 0 0 3
233 138
233 137
235 137
1 3 44 0 0 0 0 42 43 0 0 3
235 137
235 138
233 138
0 1 16 0 0 0 0 0 43 78 0 4
141 130
176 130
176 129
184 129
3 2 45 0 0 8320 0 44 47 0 0 4
341 100
357 100
357 72
380 72
2 1 46 0 0 4224 0 45 44 0 0 2
271 91
295 91
0 2 17 0 0 0 0 0 44 80 0 2
79 109
295 109
3 1 47 0 0 4224 0 46 45 0 0 2
231 91
235 91
0 2 15 0 0 0 0 0 46 77 0 2
172 100
182 100
0 1 10 0 0 0 0 0 46 79 0 2
113 82
182 82
0 1 16 0 0 4096 0 0 47 78 0 2
141 54
380 54
1 0 15 0 0 4224 0 1 0 0 0 6
172 50
172 474
171 474
171 482
172 482
172 765
1 0 16 0 0 4224 0 2 0 0 0 4
141 51
141 473
140 473
140 766
1 0 10 0 0 8320 0 3 0 0 0 4
112 51
113 51
113 765
112 765
1 0 17 0 0 12416 0 4 0 0 0 4
79 51
79 253
78 253
78 767
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
51 21 80 45
61 29 69 45
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
84 21 113 45
94 29 102 45
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
117 21 146 45
127 29 135 45
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
145 22 174 46
155 30 163 46
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
386 73 415 97
396 81 404 97
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
385 155 414 179
395 163 403 179
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
386 221 415 245
396 229 404 245
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
385 319 414 343
395 327 403 343
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
382 477 411 501
392 485 400 501
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
382 565 411 589
392 573 400 589
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
395 754 424 778
405 762 413 778
1 7
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
