CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
174 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
342 176 455 273
42991634 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 370 34 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 20592 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43485.4 0
0
13 Logic Switch~
5 261 31 0 1 11
0 9
0
0 0 20592 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43485.4 0
0
13 Logic Switch~
5 155 36 0 1 11
0 7
0
0 0 20592 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43485.4 0
0
13 Logic Switch~
5 54 36 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 20592 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
43485.4 0
0
8 2-In OR~
219 618 673 0 3 22
0 4 15 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
8157 0 0
2
43485.4 0
0
8 2-In OR~
219 539 664 0 3 22
0 6 5 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
5572 0 0
2
43485.4 0
0
6 74136~
219 471 690 0 3 22
0 7 9 5
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8901 0 0
2
43485.4 0
0
9 2-In AND~
219 474 643 0 3 22
0 9 8 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
7361 0 0
2
43485.4 0
0
8 2-In OR~
219 611 560 0 3 22
0 12 11 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
4747 0 0
2
43485.4 0
0
9 2-In AND~
219 543 594 0 3 22
0 13 7 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
972 0 0
2
43485.4 0
0
8 2-In OR~
219 466 585 0 3 22
0 14 8 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
3472 0 0
2
43485.4 0
0
8 2-In OR~
219 523 538 0 3 22
0 16 15 12
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
9998 0 0
2
43485.4 0
0
9 2-In AND~
219 472 529 0 3 22
0 14 8 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3536 0 0
2
43485.4 0
0
9 2-In AND~
219 540 484 0 3 22
0 18 8 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
4597 0 0
2
43485.4 0
0
8 2-In OR~
219 461 475 0 3 22
0 25 9 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3835 0 0
2
43485.4 0
0
8 2-In OR~
219 671 352 0 3 22
0 21 20 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3670 0 0
2
43485.4 0
0
5 7415~
219 468 426 0 4 22
0 7 14 23 22
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 7 0
1 U
5616 0 0
2
43485.4 0
0
8 2-In OR~
219 538 386 0 3 22
0 24 22 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9323 0 0
2
43485.4 0
0
9 2-In AND~
219 465 377 0 3 22
0 9 8 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
317 0 0
2
43485.4 0
0
9 2-In AND~
219 613 342 0 3 22
0 26 25 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3108 0 0
2
43485.4 0
0
8 2-In OR~
219 541 322 0 3 22
0 27 8 26
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4299 0 0
2
43485.4 0
0
8 2-In OR~
219 460 311 0 3 22
0 15 9 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9672 0 0
2
43485.4 0
0
8 2-In OR~
219 543 268 0 3 22
0 29 23 28
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7876 0 0
2
43485.4 0
0
8 2-In OR~
219 465 251 0 3 22
0 7 14 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
6369 0 0
2
43485.4 0
0
8 2-In OR~
219 596 210 0 3 22
0 31 25 30
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9172 0 0
2
43485.4 0
0
9 Inverter~
13 542 201 0 2 22
0 32 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
7100 0 0
2
43485.4 0
0
9 2-In XOR~
219 467 201 0 3 22
0 9 23 32
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3820 0 0
2
43485.4 0
0
7 Ground~
168 924 24 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7678 0 0
2
43485.4 0
0
9 CC 7-Seg~
183 924 109 0 17 19
10 33 30 28 19 17 10 3 37 2
1 1 1 1 0 1 1 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
961 0 0
2
43485.4 0
0
8 2-In OR~
219 649 154 0 3 22
0 34 9 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3178 0 0
2
43485.4 0
0
8 2-In OR~
219 579 132 0 3 22
0 35 15 34
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3409 0 0
2
43485.4 0
0
9 Inverter~
13 529 123 0 2 22
0 36 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3951 0 0
2
43485.4 0
0
6 74136~
219 466 123 0 3 22
0 7 23 36
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8885 0 0
2
43485.4 0
0
9 Inverter~
13 402 76 0 2 22
0 23 8
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3780 0 0
2
43485.4 0
0
9 Inverter~
13 292 77 0 2 22
0 9 14
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9265 0 0
2
43485.4 0
0
9 Inverter~
13 185 78 0 2 22
0 7 25
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9442 0 0
2
43485.4 0
0
68
7 3 3 0 0 4224 0 29 5 0 0 3
939 145
939 673
651 673
1 3 4 0 0 4224 0 5 6 0 0 2
605 664
572 664
3 2 5 0 0 8320 0 7 6 0 0 4
504 690
518 690
518 673
526 673
3 1 6 0 0 4224 0 8 6 0 0 4
495 643
518 643
518 655
526 655
0 1 7 0 0 4096 0 0 7 66 0 4
155 659
447 659
447 681
455 681
2 0 8 0 0 8208 0 8 0 0 59 3
450 652
450 648
404 648
0 1 9 0 0 4096 0 0 8 62 0 2
261 634
450 634
6 3 10 0 0 4224 0 29 9 0 0 3
933 145
933 560
644 560
3 2 11 0 0 4224 0 10 9 0 0 4
564 594
590 594
590 569
598 569
3 1 12 0 0 4224 0 12 9 0 0 4
556 538
590 538
590 551
598 551
0 2 7 0 0 4096 0 0 10 66 0 4
155 617
506 617
506 603
519 603
3 1 13 0 0 4224 0 11 10 0 0 2
499 585
519 585
2 0 8 0 0 4096 0 11 0 0 59 2
453 594
404 594
1 0 14 0 0 4096 0 11 0 0 0 2
453 576
295 576
2 0 15 0 0 12288 0 12 0 0 67 4
510 547
497 547
497 553
54 553
1 3 16 0 0 4224 0 12 13 0 0 2
510 529
493 529
2 0 8 0 0 0 0 13 0 0 59 2
448 538
404 538
1 0 14 0 0 0 0 13 0 0 64 2
448 520
295 520
5 3 17 0 0 8320 0 29 14 0 0 3
927 145
927 484
561 484
0 2 8 0 0 4096 0 0 14 59 0 4
404 500
508 500
508 493
516 493
3 1 18 0 0 4224 0 15 14 0 0 2
494 475
516 475
2 0 9 0 0 0 0 15 0 0 62 2
448 484
261 484
3 4 19 0 0 4224 0 16 29 0 0 3
704 352
921 352
921 145
3 2 20 0 0 4224 0 18 16 0 0 4
571 386
653 386
653 361
658 361
3 1 21 0 0 4224 0 20 16 0 0 4
634 342
653 342
653 343
658 343
4 2 22 0 0 8320 0 17 18 0 0 4
489 426
517 426
517 395
525 395
3 0 23 0 0 4096 0 17 0 0 63 2
444 435
370 435
2 0 14 0 0 0 0 17 0 0 64 2
444 426
295 426
1 0 7 0 0 0 0 17 0 0 66 2
444 417
155 417
1 3 24 0 0 4224 0 18 19 0 0 2
525 377
486 377
2 0 8 0 0 0 0 19 0 0 59 2
441 386
404 386
1 0 9 0 0 0 0 19 0 0 62 2
441 368
261 368
2 0 25 0 0 4224 0 20 0 0 65 2
589 351
193 351
1 3 26 0 0 8320 0 20 21 0 0 4
589 333
581 333
581 322
574 322
2 0 8 0 0 0 0 21 0 0 59 4
528 331
497 331
497 332
404 332
3 1 27 0 0 12416 0 22 21 0 0 4
493 311
508 311
508 313
528 313
2 0 9 0 0 0 0 22 0 0 62 2
447 320
261 320
1 0 15 0 0 0 0 22 0 0 67 2
447 302
54 302
3 3 28 0 0 4224 0 23 29 0 0 3
576 268
915 268
915 145
2 0 23 0 0 4096 0 23 0 0 63 2
530 277
370 277
1 3 29 0 0 4224 0 23 24 0 0 4
530 259
513 259
513 251
498 251
2 0 14 0 0 0 0 24 0 0 64 2
452 260
295 260
1 0 7 0 0 0 0 24 0 0 66 2
452 242
155 242
2 3 30 0 0 8320 0 29 25 0 0 3
909 145
909 210
629 210
2 0 25 0 0 0 0 25 0 0 65 4
583 219
203 219
203 220
193 220
1 2 31 0 0 4224 0 25 26 0 0 2
583 201
563 201
3 1 32 0 0 4224 0 27 26 0 0 2
500 201
527 201
2 0 23 0 0 0 0 27 0 0 63 4
451 210
375 210
375 211
370 211
1 0 9 0 0 4096 0 27 0 0 62 2
451 192
261 192
9 1 2 0 0 4224 0 29 28 0 0 2
924 67
924 32
3 1 33 0 0 4224 0 30 29 0 0 3
682 154
903 154
903 145
2 0 9 0 0 4096 0 30 0 0 62 2
636 163
261 163
3 1 34 0 0 4224 0 31 30 0 0 4
612 132
628 132
628 145
636 145
2 0 15 0 0 4096 0 31 0 0 67 2
566 141
54 141
2 1 35 0 0 4224 0 32 31 0 0 2
550 123
566 123
1 3 36 0 0 4224 0 32 33 0 0 2
514 123
499 123
2 0 23 0 0 0 0 33 0 0 63 2
450 132
370 132
1 0 7 0 0 0 0 33 0 0 66 2
450 114
155 114
2 0 8 0 0 8320 0 34 0 0 0 3
405 94
404 94
404 651
1 1 23 0 0 0 0 1 34 0 0 4
370 46
370 50
405 50
405 58
1 1 9 0 0 0 0 2 35 0 0 4
261 43
261 51
295 51
295 59
1 2 9 0 0 4224 0 2 7 0 0 5
261 43
261 676
442 676
442 699
455 699
1 0 23 0 0 4224 0 1 0 0 0 2
370 46
370 436
2 0 14 0 0 4224 0 35 0 0 14 2
295 95
295 576
2 1 25 0 0 0 0 36 15 0 0 4
188 96
193 96
193 466
448 466
1 0 7 0 0 4224 0 3 0 0 0 2
155 48
155 659
1 2 15 0 0 4224 0 4 5 0 0 5
54 48
54 733
597 733
597 682
605 682
1 1 7 0 0 0 0 3 36 0 0 4
155 48
155 52
188 52
188 60
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
354 -5 383 19
364 3 372 19
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
244 -6 273 18
254 2 262 18
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
140 -5 169 19
150 3 158 19
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
39 -5 68 19
49 3 57 19
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
