CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 35 78 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43486.4 0
0
13 Logic Switch~
5 75 80 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-7 -31 7 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
43486.4 1
0
13 Logic Switch~
5 116 80 0 1 11
0 3
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
43486.4 2
0
13 Logic Switch~
5 156 81 0 1 11
0 27
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43486.4 3
0
7 Ground~
168 534 61 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
43486.4 4
0
9 CC 7-Seg~
183 615 97 0 17 19
10 12 11 10 9 8 7 6 36 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5572 0 0
2
43486.4 5
0
8 2-In OR~
219 388 1079 0 3 22
0 13 5 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
8901 0 0
2
43486.4 6
0
8 2-In OR~
219 284 1062 0 3 22
0 15 14 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
7361 0 0
2
43486.4 7
0
6 74136~
219 211 1098 0 3 22
0 3 4 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4747 0 0
2
43486.4 8
0
9 2-In AND~
219 221 1034 0 3 22
0 16 3 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
972 0 0
2
43486.4 9
0
8 2-In OR~
219 388 901 0 3 22
0 18 17 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3472 0 0
2
43486.4 10
0
9 2-In AND~
219 303 932 0 3 22
0 4 19 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
9998 0 0
2
43486.4 11
0
8 2-In OR~
219 213 945 0 3 22
0 16 20 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3536 0 0
2
43486.4 12
0
8 2-In OR~
219 296 877 0 3 22
0 21 5 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4597 0 0
2
43486.4 13
0
9 2-In AND~
219 224 851 0 3 22
0 16 20 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3835 0 0
2
43486.4 14
0
9 2-In AND~
219 408 744 0 3 22
0 16 22 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3670 0 0
2
43486.4 15
0
8 2-In OR~
219 216 760 0 3 22
0 3 23 22
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
5616 0 0
2
43486.4 16
0
8 3-In OR~
219 401 606 0 4 22
0 26 25 24 9
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
9323 0 0
2
43486.4 17
0
5 7415~
219 342 659 0 4 22
0 27 20 4 24
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
317 0 0
2
43486.4 18
0
9 2-In AND~
219 343 606 0 3 22
0 16 3 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3108 0 0
2
43486.4 19
0
9 2-In AND~
219 344 553 0 3 22
0 28 23 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4299 0 0
2
43486.4 20
0
8 2-In OR~
219 282 530 0 3 22
0 29 16 28
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9672 0 0
2
43486.4 21
0
8 2-In OR~
219 219 511 0 3 22
0 3 5 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7876 0 0
2
43486.4 22
0
8 2-In OR~
219 406 423 0 3 22
0 30 27 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6369 0 0
2
43486.4 23
0
8 2-In OR~
219 222 402 0 3 22
0 20 4 30
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9172 0 0
2
43486.4 24
0
8 2-In OR~
219 409 299 0 3 22
0 31 23 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7100 0 0
2
43486.4 25
0
9 Inverter~
13 291 290 0 2 22
0 32 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3820 0 0
2
43486.4 26
0
6 74136~
219 229 290 0 3 22
0 27 3 32
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7678 0 0
2
43486.4 27
0
8 2-In OR~
219 408 147 0 3 22
0 3 33 12
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
961 0 0
2
43486.4 28
0
8 2-In OR~
219 311 180 0 3 22
0 34 5 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3178 0 0
2
43486.4 29
0
9 Inverter~
13 273 166 0 2 22
0 35 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3409 0 0
2
43486.4 30
0
6 74136~
219 220 166 0 3 22
0 27 4 35
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
43486.4 31
0
9 Inverter~
13 175 121 0 2 22
0 27 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8885 0 0
2
43486.4 32
0
9 Inverter~
13 132 121 0 2 22
0 3 20
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3780 0 0
2
43486.4 33
0
9 Inverter~
13 89 121 0 2 22
0 4 23
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9265 0 0
2
43486.4 34
0
63
1 0 3 0 0 4096 0 29 0 0 55 4
395 138
192 138
192 142
117 142
2 0 4 0 0 4096 0 32 0 0 50 2
204 175
75 175
2 0 5 0 0 4096 0 30 0 0 47 2
298 189
35 189
9 1 2 0 0 8320 0 6 5 0 0 4
615 55
615 47
534 47
534 55
7 3 6 0 0 4224 0 6 7 0 0 3
630 133
630 1079
421 1079
6 3 7 0 0 4224 0 6 11 0 0 3
624 133
624 901
421 901
5 3 8 0 0 4224 0 6 16 0 0 3
618 133
618 744
429 744
4 4 9 0 0 4224 0 6 18 0 0 3
612 133
612 606
434 606
3 3 10 0 0 4224 0 6 24 0 0 3
606 133
606 423
439 423
2 3 11 0 0 4224 0 6 26 0 0 3
600 133
600 299
442 299
1 3 12 0 0 8320 0 6 29 0 0 3
594 133
594 147
441 147
0 2 5 0 0 8192 0 0 7 26 0 5
37 886
37 1125
325 1125
325 1088
375 1088
1 3 13 0 0 4224 0 7 8 0 0 4
375 1070
325 1070
325 1062
317 1062
2 3 14 0 0 8320 0 8 9 0 0 4
271 1071
252 1071
252 1098
244 1098
1 3 15 0 0 4224 0 8 10 0 0 4
271 1053
250 1053
250 1034
242 1034
1 0 3 0 0 0 0 9 0 0 19 3
195 1089
119 1089
119 1043
0 2 4 0 0 4096 0 0 9 23 0 3
76 923
76 1107
195 1107
1 0 16 0 0 8192 0 10 0 0 25 3
197 1025
179 1025
179 936
2 0 3 0 0 8320 0 10 0 0 32 3
197 1043
119 1043
119 751
2 3 17 0 0 4224 0 11 12 0 0 4
375 910
337 910
337 932
324 932
1 3 18 0 0 4224 0 11 14 0 0 4
375 892
337 892
337 877
329 877
2 3 19 0 0 4224 0 12 13 0 0 4
279 941
254 941
254 945
246 945
1 0 4 0 0 8192 0 12 0 0 39 4
279 923
75 923
75 667
76 667
2 0 20 0 0 8192 0 13 0 0 29 3
200 954
135 954
135 859
1 0 16 0 0 8192 0 13 0 0 28 3
200 936
178 936
178 837
0 2 5 0 0 4096 0 0 14 47 0 3
37 520
37 886
283 886
1 3 21 0 0 4224 0 14 15 0 0 4
283 868
253 868
253 851
245 851
1 0 16 0 0 8192 0 15 0 0 30 3
200 842
178 842
178 735
0 2 20 0 0 8192 0 0 15 38 0 4
136 659
135 659
135 860
200 860
1 0 16 0 0 4096 0 16 0 0 40 3
384 735
178 735
178 597
2 3 22 0 0 8320 0 16 17 0 0 3
384 753
384 760
249 760
1 0 3 0 0 0 0 17 0 0 41 4
203 751
119 751
119 615
118 615
2 0 23 0 0 8192 0 17 0 0 42 3
203 769
93 769
93 562
3 4 24 0 0 8320 0 18 19 0 0 4
388 615
371 615
371 659
363 659
2 3 25 0 0 4224 0 18 20 0 0 2
389 606
364 606
1 3 26 0 0 8320 0 18 21 0 0 4
388 597
373 597
373 553
365 553
1 0 27 0 0 8192 0 19 0 0 48 3
318 650
156 650
156 432
0 2 20 0 0 4224 0 0 19 51 0 3
136 393
136 659
318 659
0 3 4 0 0 4096 0 0 19 50 0 3
76 411
76 668
318 668
1 0 16 0 0 0 0 20 0 0 44 3
319 597
178 597
178 539
0 2 3 0 0 0 0 0 20 46 0 3
118 502
118 615
319 615
2 0 23 0 0 8192 0 21 0 0 53 3
320 562
92 562
92 313
1 3 28 0 0 4224 0 21 22 0 0 3
320 544
320 530
315 530
2 2 16 0 0 8320 0 22 33 0 0 3
269 539
178 539
178 139
1 3 29 0 0 8320 0 22 23 0 0 4
269 521
260 521
260 511
252 511
1 0 3 0 0 0 0 23 0 0 55 3
206 502
117 502
117 299
1 2 5 0 0 4224 0 1 23 0 0 3
35 90
35 520
206 520
2 0 27 0 0 4224 0 24 0 0 56 3
393 432
156 432
156 281
1 3 30 0 0 4224 0 24 25 0 0 4
393 414
263 414
263 402
255 402
2 0 4 0 0 8320 0 25 0 0 61 3
209 411
75 411
75 98
1 2 20 0 0 0 0 25 34 0 0 3
209 393
135 393
135 139
2 1 31 0 0 4224 0 27 26 0 0 2
312 290
396 290
2 2 23 0 0 4224 0 26 35 0 0 5
396 308
92 308
92 313
92 313
92 139
1 3 32 0 0 4224 0 27 28 0 0 2
276 290
262 290
2 0 3 0 0 0 0 28 0 0 62 3
213 299
117 299
117 98
1 0 27 0 0 0 0 28 0 0 60 3
213 281
156 281
156 156
2 3 33 0 0 4224 0 29 30 0 0 4
395 156
349 156
349 180
344 180
1 2 34 0 0 4224 0 30 31 0 0 3
298 171
298 166
294 166
1 3 35 0 0 4224 0 31 32 0 0 2
258 166
253 166
1 0 27 0 0 0 0 32 0 0 63 3
204 157
156 157
156 99
1 1 4 0 0 0 0 35 2 0 0 4
92 103
92 98
75 98
75 92
1 1 3 0 0 0 0 34 3 0 0 4
135 103
135 98
116 98
116 92
1 1 27 0 0 0 0 33 4 0 0 4
178 103
178 99
156 99
156 93
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
420 856 498 871
434 867 483 878
7 GROUP F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
429 712 507 727
443 723 492 734
7 GROUP E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
438 564 515 588
448 572 504 588
7 GROUP D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
430 385 507 409
440 393 496 409
7 GROUP C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
436 262 513 286
446 270 502 286
7 GROUP B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
438 107 515 131
448 115 504 131
7 GROUP A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
144 23 169 47
152 31 160 47
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
102 22 131 46
112 30 120 46
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
62 23 87 47
70 31 78 47
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
21 22 50 46
31 30 39 46
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
