CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
110100498 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 218 57 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3932 0 0
2
43486.4 0
0
13 Logic Switch~
5 158 57 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5288 0 0
2
43486.4 1
0
13 Logic Switch~
5 38 59 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4934 0 0
2
43486.4 2
0
13 Logic Switch~
5 97 59 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5987 0 0
2
43486.4 3
0
7 Ground~
168 869 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7737 0 0
2
43486.4 0
0
9 CC 7-Seg~
183 767 354 0 18 19
10 28 25 4 20 3 14 8 2 31
1 1 1 1 0 1 1 0 2
0
0 0 21088 0
8 YELLOWCC
6 -41 62 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
4200 0 0
2
43486.4 0
0
8 3-In OR~
219 381 655 0 4 22
0 11 10 9 8
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 7 0
1 U
5780 0 0
2
43486.4 5
0
9 2-In AND~
219 302 655 0 3 22
0 13 12 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
6490 0 0
2
43486.4 6
0
9 2-In XOR~
219 297 608 0 3 22
0 12 7 11
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8663 0 0
2
43486.4 7
0
8 3-In OR~
219 439 550 0 4 22
0 16 15 9 14
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 7 0
1 U
318 0 0
2
43486.4 9
0
9 2-In AND~
219 379 549 0 3 22
0 13 17 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
348 0 0
2
43486.4 10
0
9 2-In AND~
219 375 500 0 3 22
0 18 7 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
8551 0 0
2
43486.4 11
0
8 2-In OR~
219 293 490 0 3 22
0 13 17 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7295 0 0
2
43486.4 12
0
9 2-In AND~
219 378 453 0 3 22
0 19 13 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9900 0 0
2
43486.4 14
0
8 2-In OR~
219 292 444 0 3 22
0 12 5 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
8725 0 0
2
43486.4 15
0
8 3-In OR~
219 440 354 0 4 22
0 23 22 21 20
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
366 0 0
2
43486.4 17
0
5 7415~
219 378 401 0 4 22
0 6 17 7 21
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
5762 0 0
2
43486.4 18
0
9 2-In AND~
219 379 354 0 3 22
0 13 12 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
4943 0 0
2
43486.4 19
0
9 2-In AND~
219 380 305 0 3 22
0 24 5 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3435 0 0
2
43486.4 20
0
8 3-In OR~
219 293 295 0 4 22
0 13 12 9 24
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 3 0
1 U
8705 0 0
2
43486.4 21
0
8 3-In OR~
219 293 249 0 4 22
0 7 17 6 4
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 3 0
1 U
4331 0 0
2
43486.4 23
0
8 2-In OR~
219 416 200 0 3 22
0 26 5 25
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
787 0 0
2
43486.4 25
0
9 Inverter~
13 361 191 0 2 22
0 27 26
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3655 0 0
2
43486.4 26
0
9 2-In XOR~
219 297 190 0 3 22
0 6 12 27
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6682 0 0
2
43486.4 27
0
8 3-In OR~
219 435 139 0 4 22
0 29 12 9 28
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
582 0 0
2
43486.4 29
0
9 Inverter~
13 377 130 0 2 22
0 30 29
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3125 0 0
2
43486.4 30
0
9 2-In XOR~
219 296 130 0 3 22
0 6 7 30
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5466 0 0
2
43486.4 31
0
9 Inverter~
13 237 93 0 2 22
0 6 13
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
52 0 0
2
43486.4 32
0
9 Inverter~
13 177 92 0 2 22
0 12 17
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3898 0 0
2
43486.4 33
0
9 Inverter~
13 117 93 0 2 22
0 7 5
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9413 0 0
2
43486.4 34
0
64
8 1 2 0 0 8320 0 6 5 0 0 4
788 390
788 424
869 424
869 435
0 5 3 0 0 4224 0 0 6 23 0 3
502 451
770 451
770 390
0 3 4 0 0 8192 0 0 6 43 0 5
509 249
661 249
661 425
758 425
758 390
2 0 5 0 0 4096 0 19 0 0 26 2
356 314
120 314
3 0 6 0 0 4096 0 21 0 0 36 2
280 258
218 258
2 0 5 0 0 4096 0 22 0 0 26 2
403 209
120 209
1 0 6 0 0 4096 0 24 0 0 36 2
281 181
218 181
1 0 6 0 0 0 0 27 0 0 36 2
280 121
218 121
2 0 7 0 0 4096 0 12 0 0 63 2
351 509
97 509
4 7 8 0 0 4224 0 7 6 0 0 3
414 655
782 655
782 390
3 0 9 0 0 12288 0 7 0 0 64 5
368 664
350 664
350 695
38 695
38 573
3 2 10 0 0 4224 0 8 7 0 0 2
323 655
369 655
3 1 11 0 0 8320 0 9 7 0 0 4
330 608
352 608
352 646
368 646
2 0 12 0 0 4096 0 8 0 0 61 3
278 664
158 664
158 599
1 0 13 0 0 8192 0 8 0 0 30 3
278 646
240 646
240 539
4 6 14 0 0 8320 0 10 6 0 0 4
472 550
472 552
776 552
776 390
3 2 15 0 0 8320 0 11 10 0 0 3
400 549
400 550
427 550
3 1 16 0 0 8320 0 12 10 0 0 4
396 500
409 500
409 541
426 541
2 0 17 0 0 4096 0 11 0 0 21 3
355 558
181 558
181 499
3 1 18 0 0 8320 0 13 12 0 0 3
326 490
326 491
351 491
2 0 17 0 0 0 0 13 0 0 29 2
280 499
180 499
1 0 13 0 0 0 0 13 0 0 30 2
280 481
240 481
3 0 3 0 0 128 0 14 0 0 0 3
399 453
399 451
509 451
2 0 13 0 0 4096 0 14 0 0 30 2
354 462
240 462
1 3 19 0 0 4224 0 14 15 0 0 2
354 444
325 444
2 2 5 0 0 8320 0 15 30 0 0 3
279 453
120 453
120 111
1 0 12 0 0 4096 0 15 0 0 61 2
279 435
158 435
4 4 20 0 0 8320 0 16 6 0 0 6
473 354
473 353
650 353
650 442
764 442
764 390
0 0 17 0 0 0 0 0 0 35 0 2
180 401
180 513
0 1 13 0 0 4096 0 0 11 47 0 3
240 381
240 540
355 540
3 4 21 0 0 8320 0 16 17 0 0 4
427 363
412 363
412 401
399 401
2 3 22 0 0 4224 0 16 18 0 0 2
428 354
400 354
3 1 23 0 0 8320 0 19 16 0 0 4
401 305
411 305
411 345
427 345
3 0 7 0 0 4096 0 17 0 0 63 2
354 410
97 410
2 0 17 0 0 0 0 17 0 0 58 2
354 401
180 401
1 1 6 0 0 8320 0 17 1 0 0 3
354 392
218 392
218 69
2 0 12 0 0 4096 0 18 0 0 61 2
355 363
158 363
1 0 13 0 0 0 0 18 0 0 47 2
355 345
240 345
4 1 24 0 0 8320 0 20 19 0 0 3
326 295
326 296
356 296
3 0 9 0 0 0 0 20 0 0 64 2
280 304
38 304
2 0 12 0 0 0 0 20 0 0 61 2
281 295
158 295
1 0 13 0 0 0 0 20 0 0 47 2
280 286
240 286
4 0 4 0 0 4224 0 21 0 0 0 3
326 249
509 249
509 245
2 0 17 0 0 0 0 21 0 0 58 2
281 249
180 249
1 0 7 0 0 0 0 21 0 0 63 2
280 240
97 240
3 2 25 0 0 4224 0 22 6 0 0 5
449 200
674 200
674 412
752 412
752 390
0 0 13 0 0 4224 0 0 0 57 0 2
240 188
240 406
2 1 26 0 0 4224 0 23 22 0 0 2
382 191
403 191
3 1 27 0 0 8320 0 24 23 0 0 3
330 190
330 191
346 191
2 0 12 0 0 0 0 24 0 0 61 2
281 199
158 199
4 1 28 0 0 12416 0 25 6 0 0 6
468 139
468 141
695 141
695 404
746 404
746 390
3 0 9 0 0 12288 0 25 0 0 64 4
422 148
412 148
412 159
38 159
2 0 12 0 0 12288 0 25 0 0 61 4
423 139
396 139
396 148
158 148
2 1 29 0 0 4224 0 26 25 0 0 2
398 130
422 130
3 1 30 0 0 4224 0 27 26 0 0 2
329 130
362 130
2 0 7 0 0 0 0 27 0 0 63 2
280 139
97 139
2 0 13 0 0 0 0 28 0 0 0 2
240 111
240 213
2 0 17 0 0 4224 0 29 0 0 0 2
180 110
180 409
1 1 6 0 0 0 0 28 1 0 0 3
240 75
240 69
218 69
1 1 12 0 0 0 0 29 2 0 0 3
180 74
180 69
158 69
1 1 12 0 0 4224 0 2 9 0 0 3
158 69
158 599
281 599
1 1 7 0 0 0 0 30 4 0 0 3
120 75
120 71
97 71
1 2 7 0 0 4224 0 4 9 0 0 3
97 71
97 617
281 617
1 3 9 0 0 4224 0 3 10 0 0 5
38 71
38 574
409 574
409 559
426 559
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
521 621 548 643
530 628 538 644
1 G
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
522 517 549 539
531 525 539 541
1 F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
524 415 551 437
533 422 541 438
1 E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
525 317 548 339
532 325 540 341
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
523 213 546 235
530 220 538 236
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
523 171 546 193
530 178 538 194
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
525 108 548 130
532 115 540 131
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
202 0 231 24
212 8 220 24
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
141 0 166 24
149 8 157 24
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
80 0 109 24
90 8 98 24
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
25 0 50 24
33 8 41 24
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
