CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 331 27 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -27 8 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3701 0 0
2
43484.8 0
0
13 Logic Switch~
5 242 28 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -28 8 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6316 0 0
2
43484.8 0
0
13 Logic Switch~
5 151 27 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8734 0 0
2
43484.8 0
0
13 Logic Switch~
5 63 29 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7988 0 0
2
43484.8 0
0
7 Ground~
168 935 41 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3217 0 0
2
43484.9 0
0
8 2-In OR~
219 576 751 0 3 22
0 6 5 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3965 0 0
2
43484.9 0
0
8 2-In OR~
219 508 704 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
8239 0 0
2
43484.9 0
0
6 74136~
219 441 737 0 3 22
0 10 9 7
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
828 0 0
2
43484.8 0
0
9 2-In AND~
219 447 686 0 3 22
0 9 3 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
6187 0 0
2
43484.8 0
0
8 2-In OR~
219 581 599 0 3 22
0 13 12 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
7107 0 0
2
43484.8 0
0
9 2-In AND~
219 519 636 0 3 22
0 14 10 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
6433 0 0
2
43484.8 0
0
8 2-In OR~
219 440 612 0 3 22
0 15 3 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
8559 0 0
2
43484.8 0
0
8 2-In OR~
219 507 572 0 3 22
0 16 5 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3674 0 0
2
43484.8 0
0
9 2-In AND~
219 448 543 0 3 22
0 15 3 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
5697 0 0
2
43484.8 0
0
9 2-In AND~
219 523 504 0 3 22
0 18 3 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3805 0 0
2
43484.8 0
0
8 2-In OR~
219 441 471 0 3 22
0 19 9 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
5219 0 0
2
43484.8 0
0
8 2-In OR~
219 689 361 0 3 22
0 22 21 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3795 0 0
2
43484.8 0
0
9 2-In AND~
219 617 334 0 3 22
0 23 19 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3637 0 0
2
43484.8 0
0
8 2-In OR~
219 556 393 0 3 22
0 25 24 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3226 0 0
2
43484.8 0
0
5 7415~
219 495 421 0 4 22
0 10 15 26 24
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
6966 0 0
2
43484.8 0
0
9 2-In AND~
219 495 369 0 3 22
0 9 3 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9796 0 0
2
43484.8 0
0
8 2-In OR~
219 514 316 0 3 22
0 27 3 23
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5952 0 0
2
43484.8 0
0
8 2-In OR~
219 447 293 0 3 22
0 5 9 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3649 0 0
2
43484.8 0
0
8 2-In OR~
219 517 247 0 3 22
0 29 26 28
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3716 0 0
2
43484.8 0
0
8 2-In OR~
219 447 231 0 3 22
0 10 15 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
4797 0 0
2
43484.8 0
0
8 2-In OR~
219 517 184 0 3 22
0 31 19 30
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4681 0 0
2
43484.8 0
0
6 74136~
219 450 169 0 3 22
0 9 3 31
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9730 0 0
2
43484.8 0
0
8 2-In OR~
219 614 131 0 3 22
0 33 9 32
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9874 0 0
2
43484.8 0
0
8 2-In OR~
219 552 106 0 3 22
0 34 5 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
364 0 0
2
43484.8 0
0
9 Inverter~
13 497 89 0 2 22
0 35 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3656 0 0
2
43484.8 0
0
6 74136~
219 453 89 0 3 22
0 10 26 35
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3131 0 0
2
43484.8 0
0
9 Inverter~
13 372 57 0 2 22
0 26 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6772 0 0
2
43484.8 0
0
9 Inverter~
13 280 60 0 2 22
0 9 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9557 0 0
2
43484.8 0
0
9 Inverter~
13 183 60 0 2 22
0 10 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
5789 0 0
2
43484.8 0
0
9 Inverter~
13 92 61 0 2 22
0 5 36
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7328 0 0
2
43484.8 0
0
9 CC 7-Seg~
183 935 119 0 17 19
10 32 30 28 20 17 11 4 37 2
1 1 1 1 0 1 1 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
4799 0 0
2
43484.8 0
0
72
0 2 3 0 0 4096 0 0 21 61 0 2
393 378
471 378
0 2 3 0 0 0 0 0 27 61 0 2
393 178
434 178
1 9 2 0 0 4224 0 5 36 0 0 2
935 49
935 77
3 7 4 0 0 8320 0 6 36 0 0 3
609 751
950 751
950 155
0 2 5 0 0 4096 0 0 6 72 0 2
63 760
563 760
3 1 6 0 0 8320 0 7 6 0 0 4
541 704
555 704
555 742
563 742
3 2 7 0 0 8320 0 8 7 0 0 4
474 737
487 737
487 713
495 713
3 1 8 0 0 4224 0 9 7 0 0 4
468 686
487 686
487 695
495 695
0 2 9 0 0 4096 0 0 8 66 0 2
242 746
425 746
0 1 10 0 0 4096 0 0 8 69 0 2
151 728
425 728
0 2 3 0 0 0 0 0 9 61 0 2
393 695
423 695
0 1 9 0 0 0 0 0 9 66 0 2
242 677
423 677
3 6 11 0 0 8320 0 10 36 0 0 3
614 599
944 599
944 155
3 2 12 0 0 8320 0 11 10 0 0 4
540 636
560 636
560 608
568 608
3 1 13 0 0 4224 0 13 10 0 0 4
540 572
560 572
560 590
568 590
0 2 10 0 0 4096 0 0 11 69 0 2
151 645
495 645
3 1 14 0 0 8320 0 12 11 0 0 4
473 612
487 612
487 627
495 627
0 2 3 0 0 0 0 0 12 61 0 2
393 621
427 621
0 1 15 0 0 4096 0 0 12 64 0 2
301 603
427 603
0 2 5 0 0 0 0 0 13 72 0 2
63 581
494 581
3 1 16 0 0 8320 0 14 13 0 0 4
469 543
486 543
486 563
494 563
0 2 3 0 0 0 0 0 14 61 0 2
393 552
424 552
0 1 15 0 0 0 0 0 14 64 0 2
301 534
424 534
3 5 17 0 0 4224 0 15 36 0 0 3
544 504
938 504
938 155
0 2 3 0 0 4096 0 0 15 61 0 2
393 513
499 513
3 1 18 0 0 8320 0 16 15 0 0 4
474 471
491 471
491 495
499 495
0 2 9 0 0 4096 0 0 16 66 0 2
242 480
428 480
0 1 19 0 0 4096 0 0 16 67 0 2
204 462
428 462
3 4 20 0 0 4224 0 17 36 0 0 3
722 361
932 361
932 155
3 2 21 0 0 4224 0 19 17 0 0 4
589 393
668 393
668 370
676 370
3 1 22 0 0 4224 0 18 17 0 0 4
638 334
668 334
668 352
676 352
0 2 19 0 0 4096 0 0 18 67 0 2
204 343
593 343
3 1 23 0 0 4224 0 22 18 0 0 4
547 316
585 316
585 325
593 325
4 2 24 0 0 4224 0 20 19 0 0 4
516 421
535 421
535 402
543 402
3 1 25 0 0 4224 0 21 19 0 0 4
516 369
535 369
535 384
543 384
0 3 26 0 0 4096 0 0 20 63 0 2
331 430
471 430
0 2 15 0 0 4096 0 0 20 64 0 2
301 421
471 421
0 1 10 0 0 0 0 0 20 69 0 2
151 412
471 412
0 1 9 0 0 4096 0 0 21 66 0 2
242 360
471 360
0 2 3 0 0 4096 0 0 22 61 0 2
393 325
501 325
3 1 27 0 0 8320 0 23 22 0 0 4
480 293
493 293
493 307
501 307
0 2 9 0 0 0 0 0 23 66 0 2
242 302
434 302
0 1 5 0 0 16 0 0 23 72 0 3
63 283
434 283
434 284
3 3 28 0 0 4224 0 24 36 0 0 3
550 247
926 247
926 155
0 2 26 0 0 4096 0 0 24 63 0 2
331 256
504 256
3 1 29 0 0 4224 0 25 24 0 0 4
480 231
496 231
496 238
504 238
0 2 15 0 0 0 0 0 25 64 0 2
301 240
434 240
0 1 10 0 0 0 0 0 25 69 0 2
151 222
434 222
3 2 30 0 0 4224 0 26 36 0 0 3
550 184
920 184
920 155
0 2 19 0 0 0 0 0 26 67 0 2
204 193
504 193
3 1 31 0 0 4224 0 27 26 0 0 4
483 169
496 169
496 175
504 175
0 1 9 0 0 0 0 0 27 66 0 2
242 160
434 160
3 1 32 0 0 4224 0 28 36 0 0 5
647 131
874 131
874 158
914 158
914 155
0 2 9 0 0 4096 0 0 28 66 0 2
242 140
601 140
3 1 33 0 0 8320 0 29 28 0 0 4
585 106
593 106
593 122
601 122
0 2 5 0 0 0 0 0 29 72 0 2
63 115
539 115
2 1 34 0 0 4224 0 30 29 0 0 4
518 89
531 89
531 97
539 97
1 3 35 0 0 4224 0 30 31 0 0 2
482 89
486 89
0 2 26 0 0 0 0 0 31 63 0 2
331 98
437 98
0 1 10 0 0 0 0 0 31 69 0 2
151 80
437 80
2 0 3 0 0 4224 0 32 0 0 0 2
393 57
393 809
0 1 26 0 0 0 0 0 32 63 0 2
331 57
357 57
1 0 26 0 0 4224 0 1 0 0 0 2
331 39
331 813
2 0 15 0 0 4224 0 33 0 0 0 2
301 60
301 814
0 1 9 0 0 0 0 0 33 66 0 3
242 59
242 60
265 60
1 0 9 0 0 4224 0 2 0 0 0 2
242 40
242 813
2 0 19 0 0 4224 0 34 0 0 0 2
204 60
204 812
0 1 10 0 0 0 0 0 34 69 0 3
151 59
151 60
168 60
1 0 10 0 0 4224 0 3 0 0 0 2
151 39
151 816
2 0 36 0 0 4224 0 35 0 0 0 2
113 61
113 816
0 1 5 0 0 0 0 0 35 72 0 3
63 59
63 61
77 61
1 0 5 0 0 4224 0 4 0 0 0 2
63 41
63 817
1
-16 0 0 0 700 0 0 0 0 10 2 1 34
8 Hobo Std
0 0 0 88
990 160 1166 268
1002 169 1153 257
88 Balaba, Napthali A.
Opelinia, Prince Lonito
Hinay, Diomedes Jr.
Villorejo, Glaiza Mae
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
