CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
64 C:\Users\REY MARK\Desktop\CicMaker2000\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 260 55 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 194 56 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 125 56 0 1 11
0 17
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 52 55 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 493 768 0 3 22
0 14 13 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
8157 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 410 712 0 3 22
0 16 15 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
5572 0 0
2
5.89878e-315 0
0
6 74136~
219 332 741 0 3 22
0 17 11 15
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8901 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 339 684 0 3 22
0 11 18 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
7361 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 469 608 0 3 22
0 20 19 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
4747 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 392 636 0 3 22
0 21 17 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
972 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 328 616 0 3 22
0 22 18 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3472 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 383 578 0 3 22
0 23 13 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
9998 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 335 561 0 3 22
0 22 18 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3536 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 413 509 0 3 22
0 24 18 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4597 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 335 494 0 3 22
0 25 11 24
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3835 0 0
2
5.89878e-315 0
0
8 3-In OR~
219 558 399 0 4 22
0 28 27 26 6
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
3670 0 0
2
5.89878e-315 0
0
5 7415~
219 358 449 0 4 22
0 17 22 10 26
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
5616 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 359 407 0 3 22
0 11 18 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9323 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 465 373 0 3 22
0 29 25 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
317 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 396 355 0 3 22
0 30 18 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3108 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 328 346 0 3 22
0 13 11 30
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4299 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 413 305 0 3 22
0 31 10 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9672 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 337 295 0 3 22
0 17 22 31
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7876 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 435 252 0 3 22
0 32 25 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6369 0 0
2
5.89878e-315 0
0
9 Inverter~
13 402 221 0 2 22
0 12 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
9172 0 0
2
5.89878e-315 0
0
6 74136~
219 342 238 0 3 22
0 11 10 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7100 0 0
2
5.89878e-315 0
0
7 Ground~
168 734 66 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
5.89878e-315 0
0
9 CC 7-Seg~
183 707 149 0 17 19
10 9 8 7 6 5 4 3 36 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7678 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 465 119 0 3 22
0 11 33 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
961 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 409 175 0 3 22
0 34 13 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3178 0 0
2
5.89878e-315 0
0
9 Inverter~
13 394 127 0 2 22
0 35 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3409 0 0
2
5.89878e-315 0
0
6 74136~
219 346 149 0 3 22
0 17 10 35
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
5.89878e-315 0
0
9 Inverter~
13 295 96 0 2 22
0 10 18
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8885 0 0
2
5.89878e-315 0
0
9 Inverter~
13 219 96 0 2 22
0 11 22
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3780 0 0
2
5.89878e-315 0
0
9 Inverter~
13 149 95 0 2 22
0 17 25
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9265 0 0
2
5.89878e-315 0
0
70
7 3 3 0 0 4224 0 28 5 0 0 3
722 185
722 768
526 768
6 3 4 0 0 4224 0 28 9 0 0 3
716 185
716 608
502 608
5 3 5 0 0 4224 0 28 14 0 0 3
710 185
710 509
434 509
4 4 6 0 0 4224 0 28 16 0 0 3
704 185
704 399
591 399
3 3 7 0 0 8320 0 28 22 0 0 3
698 185
698 305
446 305
2 3 8 0 0 8320 0 28 24 0 0 3
692 185
692 252
468 252
1 9 2 0 0 8320 0 27 28 0 0 4
734 60
706 60
706 107
707 107
1 3 9 0 0 8320 0 28 29 0 0 5
686 185
686 188
506 188
506 119
498 119
2 0 10 0 0 4096 0 26 0 0 67 2
326 247
260 247
1 0 11 0 0 4096 0 26 0 0 68 2
326 229
194 229
1 3 12 0 0 8320 0 25 26 0 0 3
387 221
375 221
375 238
2 0 13 0 0 4096 0 5 0 0 70 2
480 777
52 777
3 1 14 0 0 8320 0 6 5 0 0 3
443 712
480 712
480 759
3 2 15 0 0 4224 0 7 6 0 0 3
365 741
397 741
397 721
3 1 16 0 0 4224 0 8 6 0 0 3
360 684
397 684
397 703
2 0 11 0 0 0 0 7 0 0 68 2
316 750
194 750
1 0 17 0 0 4096 0 7 0 0 69 2
316 732
125 732
2 0 18 0 0 4096 0 8 0 0 61 2
315 693
298 693
1 0 11 0 0 0 0 8 0 0 68 2
315 675
194 675
3 2 19 0 0 4224 0 10 9 0 0 3
413 636
456 636
456 617
3 1 20 0 0 4224 0 12 9 0 0 3
416 578
456 578
456 599
2 0 17 0 0 4096 0 10 0 0 69 2
368 645
125 645
1 3 21 0 0 4224 0 10 11 0 0 3
368 627
368 616
361 616
2 0 18 0 0 0 0 11 0 0 61 2
315 625
298 625
1 0 22 0 0 4096 0 11 0 0 62 2
315 607
222 607
2 0 13 0 0 0 0 12 0 0 70 2
370 587
52 587
3 1 23 0 0 4224 0 13 12 0 0 3
356 561
370 561
370 569
2 0 18 0 0 0 0 13 0 0 61 2
311 570
298 570
1 0 22 0 0 0 0 13 0 0 62 2
311 552
222 552
2 0 18 0 0 4096 0 14 0 0 61 2
389 518
298 518
3 1 24 0 0 4224 0 15 14 0 0 3
368 494
389 494
389 500
2 0 11 0 0 0 0 15 0 0 68 2
322 503
194 503
1 0 25 0 0 4096 0 15 0 0 63 2
322 485
152 485
4 3 26 0 0 4224 0 17 16 0 0 4
379 449
539 449
539 408
545 408
3 2 27 0 0 4224 0 18 16 0 0 4
380 407
528 407
528 399
546 399
3 1 28 0 0 4224 0 19 16 0 0 3
486 373
545 373
545 390
3 0 10 0 0 4096 0 17 0 0 67 2
334 458
260 458
2 0 22 0 0 4096 0 17 0 0 62 2
334 449
222 449
1 0 17 0 0 0 0 17 0 0 69 2
334 440
125 440
2 0 18 0 0 0 0 18 0 0 61 2
335 416
298 416
1 0 11 0 0 4096 0 18 0 0 68 2
335 398
194 398
2 0 25 0 0 4096 0 19 0 0 63 2
441 382
152 382
3 1 29 0 0 4224 0 20 19 0 0 3
429 355
441 355
441 364
2 0 18 0 0 0 0 20 0 0 61 2
383 364
298 364
1 3 30 0 0 4224 0 20 21 0 0 2
383 346
361 346
2 0 11 0 0 0 0 21 0 0 68 2
315 355
194 355
1 0 13 0 0 0 0 21 0 0 70 2
315 337
52 337
2 0 10 0 0 4096 0 22 0 0 67 2
400 314
260 314
1 3 31 0 0 8320 0 22 23 0 0 3
400 296
400 295
370 295
2 0 22 0 0 0 0 23 0 0 62 2
324 304
222 304
1 0 17 0 0 0 0 23 0 0 69 2
324 286
125 286
2 0 25 0 0 0 0 24 0 0 63 2
422 261
152 261
2 1 32 0 0 8320 0 25 24 0 0 3
423 221
422 221
422 243
1 0 11 0 0 4096 0 29 0 0 68 2
452 110
194 110
3 2 33 0 0 4224 0 30 29 0 0 3
442 175
442 128
452 128
2 0 13 0 0 0 0 30 0 0 70 2
396 184
52 184
2 1 34 0 0 4224 0 31 30 0 0 4
415 127
415 148
396 148
396 166
1 3 35 0 0 4224 0 31 32 0 0 2
379 127
379 149
2 0 10 0 0 0 0 32 0 0 67 2
330 158
260 158
1 0 17 0 0 0 0 32 0 0 69 2
330 140
125 140
2 0 18 0 0 4224 0 33 0 0 0 2
298 114
298 695
2 0 22 0 0 4224 0 34 0 0 0 2
222 114
222 611
2 0 25 0 0 4224 0 35 0 0 0 2
152 113
152 488
1 0 17 0 0 0 0 35 0 0 69 2
152 77
125 77
1 0 11 0 0 0 0 34 0 0 68 2
222 78
194 78
1 0 10 0 0 0 0 33 0 0 67 2
298 78
260 78
1 0 10 0 0 4224 0 1 0 0 0 2
260 67
260 461
1 0 11 0 0 4224 0 2 0 0 0 2
194 68
194 754
1 0 17 0 0 4224 0 3 0 0 0 2
125 68
125 734
1 0 13 0 0 4224 0 4 0 0 0 2
52 67
52 779
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
45 3 74 27
55 11 63 27
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
114 2 143 26
124 10 132 26
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
190 3 219 27
200 11 208 27
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
255 -1 284 23
265 7 273 23
1 D
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
