CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
38
13 Logic Switch~
5 847 87 0 1 11
0 26
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 589 86 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 366 81 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -22 8 -14
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9968 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 147 80 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9281 0 0
2
5.89878e-315 0
0
7 Ground~
168 1099 504 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8464 0 0
2
5.89878e-315 0
0
9 CC 7-Seg~
183 1099 580 0 17 19
10 9 8 7 6 5 4 3 38 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7168 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 241 509 0 3 22
0 10 11 3
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U8C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3171 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 613 578 0 3 22
0 12 13 10
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U8B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
4139 0 0
2
5.89878e-315 0
0
9 2-In XOR~
219 528 531 0 3 22
0 14 15 13
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U2C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
6435 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 961 520 0 3 22
0 16 14 12
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U7D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
5283 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 439 498 0 3 22
0 18 17 4
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U8A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
6874 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 560 363 0 3 22
0 19 15 18
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U7C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
5305 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 1025 329 0 3 22
0 16 20 19
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U6D
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
34 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 314 391 0 3 22
0 21 11 17
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U6C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
969 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 1044 225 0 3 22
0 16 20 21
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U7B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8402 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 481 274 0 3 22
0 14 23 22
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U6B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3751 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 937 344 0 3 22
0 16 22 5
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U7A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
4292 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 850 510 0 3 22
0 25 24 6
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U6A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
6118 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 883 233 0 3 22
0 26 27 25
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U5D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
34 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 662 235 0 3 22
0 20 15 27
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U5C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
6357 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 639 515 0 3 22
0 28 29 24
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U4D
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
319 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 777 508 0 3 22
0 16 14 28
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U5B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3976 0 0
2
5.89878e-315 0
0
9 2-In AND~
219 508 482 0 3 22
0 30 23 29
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7634 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 907 442 0 3 22
0 16 31 30
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U4C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
523 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 395 424 0 3 22
0 14 11 31
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U4B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6748 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 708 329 0 3 22
0 26 32 7
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U4A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6901 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 517 247 0 3 22
0 20 15 32
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U3D
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
842 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 640 408 0 3 22
0 33 23 8
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U3C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3277 0 0
2
5.89878e-315 0
0
9 Inverter~
13 777 376 0 2 22
0 34 33
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
4212 0 0
2
5.89878e-315 0
0
9 2-In XOR~
219 777 321 0 3 22
0 26 14 34
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U2B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4720 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 485 353 0 3 22
0 14 35 9
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U3B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5551 0 0
2
5.89878e-315 0
0
8 2-In OR~
219 259 303 0 3 22
0 36 11 35
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U3A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6986 0 0
2
5.89878e-315 0
0
9 Inverter~
13 922 268 0 2 22
0 37 36
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
8745 0 0
2
5.89878e-315 0
0
9 2-In XOR~
219 922 210 0 3 22
0 26 15 37
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U2A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9592 0 0
2
5.89878e-315 0
0
9 Inverter~
13 990 126 0 2 22
0 26 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8748 0 0
2
5.89878e-315 0
0
9 Inverter~
13 727 128 0 2 22
0 14 20
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
7168 0 0
2
5.89878e-315 0
0
9 Inverter~
13 470 135 0 2 22
0 15 23
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
631 0 0
2
5.89878e-315 0
0
9 Inverter~
13 202 140 0 2 22
0 11 39
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 1 1 0
1 U
9466 0 0
2
5.89878e-315 0
0
67
1 9 2 0 0 4224 0 5 6 0 0 2
1099 512
1099 538
3 7 3 0 0 8320 0 7 6 0 0 4
244 539
244 686
1114 686
1114 616
3 6 4 0 0 8320 0 11 6 0 0 4
442 528
442 675
1108 675
1108 616
3 5 5 0 0 8320 0 17 6 0 0 5
935 367
1012 367
1012 667
1102 667
1102 616
3 4 6 0 0 8320 0 18 6 0 0 4
853 540
853 659
1096 659
1096 616
3 3 7 0 0 12416 0 26 6 0 0 5
711 359
732 359
732 652
1090 652
1090 616
3 2 8 0 0 12416 0 28 6 0 0 5
643 438
719 438
719 642
1084 642
1084 616
3 1 9 0 0 8320 0 31 6 0 0 4
488 383
488 631
1078 631
1078 616
3 1 10 0 0 4224 0 8 7 0 0 4
616 608
318 608
318 493
253 493
0 2 11 0 0 4096 0 0 7 24 0 3
147 375
147 493
235 493
3 1 12 0 0 8320 0 10 8 0 0 3
959 543
959 562
625 562
3 2 13 0 0 8320 0 9 8 0 0 3
531 561
531 562
607 562
0 1 14 0 0 8192 0 0 9 16 0 3
589 480
589 512
540 512
0 2 15 0 0 4096 0 0 9 36 0 5
369 213
369 469
481 469
481 512
522 512
0 1 16 0 0 4096 0 0 10 43 0 3
993 426
993 498
968 498
0 2 14 0 0 8320 0 0 10 45 0 4
589 391
589 480
950 480
950 498
3 2 17 0 0 12416 0 14 11 0 0 4
317 421
365 421
365 482
433 482
3 1 18 0 0 8320 0 12 11 0 0 4
558 386
558 439
451 439
451 482
0 2 15 0 0 0 0 0 12 62 0 5
366 170
442 170
442 321
549 321
549 341
3 1 19 0 0 8320 0 13 12 0 0 5
1028 359
1028 397
688 397
688 341
567 341
0 1 16 0 0 8192 0 0 13 43 0 5
993 185
1016 185
1016 292
1037 292
1037 313
0 2 20 0 0 12288 0 0 13 35 0 5
730 177
823 177
823 309
1019 309
1019 313
3 1 21 0 0 8320 0 15 14 0 0 5
1042 248
1042 409
452 409
452 375
326 375
0 2 11 0 0 8192 0 0 14 59 0 3
147 287
147 375
308 375
2 1 16 0 0 0 0 35 15 0 0 3
993 144
1051 144
1051 203
0 2 20 0 0 4224 0 0 15 35 0 3
730 153
1033 153
1033 203
3 2 22 0 0 12416 0 16 17 0 0 6
484 304
545 304
545 264
909 264
909 322
926 322
0 1 14 0 0 0 0 0 16 56 0 3
589 175
493 175
493 258
0 2 23 0 0 8192 0 0 16 52 0 3
473 217
475 217
475 258
0 1 16 0 0 0 0 0 17 43 0 3
993 317
944 317
944 322
3 2 24 0 0 4224 0 21 18 0 0 4
642 545
825 545
825 494
844 494
3 1 25 0 0 4224 0 19 18 0 0 3
881 256
881 494
862 494
0 1 26 0 0 4096 0 0 19 54 0 3
847 179
890 179
890 211
3 2 27 0 0 4224 0 20 19 0 0 4
660 258
855 258
855 211
872 211
2 1 20 0 0 0 0 36 20 0 0 3
730 146
730 213
669 213
0 2 15 0 0 8192 0 0 20 62 0 3
366 191
366 213
651 213
3 1 28 0 0 4224 0 22 21 0 0 4
775 531
677 531
677 499
651 499
3 2 29 0 0 4224 0 23 21 0 0 4
506 505
616 505
616 499
633 499
0 1 16 0 0 8192 0 0 22 43 0 3
969 426
969 486
784 486
0 2 14 0 0 0 0 0 22 56 0 4
589 161
754 161
754 486
766 486
3 1 30 0 0 4224 0 24 23 0 0 4
910 472
534 472
534 460
515 460
0 2 23 0 0 8320 0 0 23 52 0 4
473 161
436 161
436 460
497 460
2 1 16 0 0 4224 0 35 24 0 0 3
993 144
993 426
919 426
3 2 31 0 0 4224 0 25 24 0 0 4
398 454
873 454
873 426
901 426
0 1 14 0 0 0 0 0 25 56 0 4
589 337
589 391
407 391
407 408
0 2 11 0 0 8320 0 0 25 59 0 4
147 120
181 120
181 408
389 408
0 1 26 0 0 4096 0 0 26 54 0 3
847 272
720 272
720 313
3 2 32 0 0 4224 0 27 26 0 0 3
520 277
702 277
702 313
2 1 20 0 0 0 0 36 27 0 0 3
730 146
529 146
529 231
0 2 15 0 0 0 0 0 27 62 0 4
366 121
456 121
456 231
511 231
2 1 33 0 0 8320 0 29 28 0 0 3
780 394
780 392
652 392
2 2 23 0 0 0 0 37 28 0 0 4
473 153
473 217
634 217
634 392
3 1 34 0 0 4224 0 30 29 0 0 2
780 351
780 358
0 1 26 0 0 4096 0 0 30 61 0 3
847 162
847 302
789 302
0 2 14 0 0 0 0 0 30 56 0 4
589 116
692 116
692 302
771 302
1 1 14 0 0 0 0 2 31 0 0 3
589 98
589 337
497 337
3 2 35 0 0 4224 0 32 31 0 0 3
262 333
479 333
479 337
2 1 36 0 0 8320 0 33 32 0 0 3
925 286
925 287
271 287
1 2 11 0 0 0 0 4 32 0 0 3
147 92
147 287
253 287
3 1 37 0 0 4224 0 34 33 0 0 2
925 240
925 250
1 1 26 0 0 0 0 1 34 0 0 4
847 99
847 163
934 163
934 191
1 2 15 0 0 8320 0 3 34 0 0 3
366 93
366 191
916 191
1 0 15 0 0 0 0 3 0 0 66 2
366 93
442 93
1 1 26 0 0 4224 0 1 35 0 0 3
847 99
993 99
993 108
1 1 14 0 0 0 0 2 36 0 0 3
589 98
730 98
730 110
1 1 15 0 0 0 0 3 37 0 0 3
366 93
473 93
473 117
1 1 11 0 0 0 0 4 38 0 0 3
147 92
205 92
205 122
11
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
487 82 523 113
497 90 512 111
1 B
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
1031 84 1068 115
1041 92 1057 113
1 D
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
473 380 509 411
484 388 497 409
1 A
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
624 433 662 464
635 441 650 462
1 B
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
693 355 730 386
704 363 718 384
1 C
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
838 536 871 567
846 544 862 565
1 D
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
916 358 954 389
927 366 942 387
1 E
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
425 525 462 556
436 533 450 554
1 F
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
225 536 264 567
236 544 252 565
1 G
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
215 83 245 114
223 91 236 112
1 A
-16 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 1
738 81 769 112
746 89 760 110
1 C
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
