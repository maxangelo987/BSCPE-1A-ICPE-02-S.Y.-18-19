CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 12 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
9437202 0
0
2 

2 

0
0
0
36
13 Logic Switch~
5 222 123 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43490.4 0
0
13 Logic Switch~
5 159 122 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
43490.4 1
0
13 Logic Switch~
5 287 121 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43490.4 2
0
13 Logic Switch~
5 92 122 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
43490.4 3
0
7 Ground~
168 846 452 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
43490.4 4
0
9 CC 7-Seg~
183 846 535 0 17 19
10 9 8 7 3 6 5 4 37 2
1 0 1 1 0 1 1 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5572 0 0
2
43490.4 5
0
8 2-In OR~
219 468 1073 0 3 22
0 15 19 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
8901 0 0
2
43490.4 6
0
8 2-In OR~
219 414 1045 0 3 22
0 16 20 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
7361 0 0
2
43490.4 7
0
9 2-In XOR~
219 354 1054 0 3 22
0 21 13 20
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4747 0 0
2
43490.4 8
0
9 2-In AND~
219 360 1005 0 3 22
0 13 12 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
972 0 0
2
43490.4 9
0
8 2-In OR~
219 469 897 0 3 22
0 23 22 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3472 0 0
2
43490.4 10
0
9 2-In AND~
219 423 934 0 3 22
0 14 21 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
9998 0 0
2
43490.4 11
0
8 2-In OR~
219 354 898 0 3 22
0 24 12 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3536 0 0
2
43490.4 12
0
8 2-In OR~
219 408 854 0 3 22
0 25 19 23
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
4597 0 0
2
43490.4 13
0
9 2-In AND~
219 368 820 0 3 22
0 24 12 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3835 0 0
2
43490.4 14
0
9 2-In AND~
219 481 751 0 3 22
0 26 12 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3670 0 0
2
43490.4 15
0
8 2-In OR~
219 356 729 0 3 22
0 13 27 26
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
5616 0 0
2
43490.4 16
0
8 3-In OR~
219 502 593 0 4 22
0 29 11 28 3
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
9323 0 0
2
43490.4 17
0
5 7415~
219 364 652 0 4 22
0 21 24 30 28
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 7 0
1 U
317 0 0
2
43490.4 18
0
9 2-In AND~
219 362 605 0 3 22
0 13 12 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3108 0 0
2
43490.4 19
0
9 2-In AND~
219 467 562 0 3 22
0 31 27 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
4299 0 0
2
43490.4 20
0
8 2-In OR~
219 402 545 0 3 22
0 10 12 31
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9672 0 0
2
43490.4 21
0
8 2-In OR~
219 353 516 0 3 22
0 19 13 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7876 0 0
2
43490.4 22
0
8 2-In OR~
219 461 455 0 3 22
0 32 30 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6369 0 0
2
43490.4 23
0
8 2-In OR~
219 353 424 0 3 22
0 21 24 32
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9172 0 0
2
43490.4 24
0
8 2-In OR~
219 459 355 0 3 22
0 33 27 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7100 0 0
2
43490.4 25
0
9 Inverter~
13 420 320 0 2 22
0 34 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3820 0 0
2
43490.4 26
0
9 2-In XOR~
219 355 320 0 3 22
0 13 30 34
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7678 0 0
2
43490.4 27
0
8 2-In OR~
219 536 253 0 3 22
0 35 13 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
961 0 0
2
43490.4 28
0
8 2-In OR~
219 473 234 0 3 22
0 17 19 35
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3178 0 0
2
43490.4 29
0
9 Inverter~
13 426 213 0 2 22
0 18 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3409 0 0
2
43490.4 30
0
6 74136~
219 354 213 0 3 22
0 21 30 18
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
43490.4 31
0
9 Inverter~
13 312 153 0 2 22
0 30 12
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8885 0 0
2
43490.4 32
0
9 Inverter~
13 246 156 0 2 22
0 13 24
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3780 0 0
2
43490.4 33
0
9 Inverter~
13 181 154 0 2 22
0 21 27
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9265 0 0
2
43490.4 34
0
9 Inverter~
13 116 154 0 2 22
0 19 36
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9442 0 0
2
43490.4 35
0
72
1 9 2 0 0 4224 0 5 6 0 0 2
846 460
846 493
4 4 3 0 0 4224 0 18 6 0 0 3
535 593
843 593
843 571
3 7 4 0 0 16512 0 7 6 0 0 5
501 1073
644 1073
644 1072
861 1072
861 571
3 6 5 0 0 4224 0 11 6 0 0 3
502 897
855 897
855 571
3 5 6 0 0 4224 0 16 6 0 0 3
502 751
849 751
849 571
3 3 7 0 0 4224 0 24 6 0 0 5
494 455
787 455
787 585
837 585
837 571
3 2 8 0 0 4224 0 26 6 0 0 5
492 355
798 355
798 577
831 577
831 571
3 1 9 0 0 8320 0 29 6 0 0 4
569 253
810 253
810 571
825 571
3 1 10 0 0 8320 0 23 22 0 0 3
386 516
389 516
389 536
2 3 11 0 0 4224 0 18 20 0 0 4
490 593
391 593
391 605
383 605
2 0 12 0 0 4096 0 10 0 0 61 2
336 1014
315 1014
1 0 13 0 0 4096 0 10 0 0 70 2
336 996
223 996
2 0 12 0 0 0 0 13 0 0 61 4
341 907
328 907
328 908
315 908
3 1 14 0 0 8320 0 13 12 0 0 3
387 898
399 898
399 925
3 1 15 0 0 8320 0 8 7 0 0 4
447 1045
448 1045
448 1064
455 1064
3 1 16 0 0 8320 0 10 8 0 0 4
381 1005
388 1005
388 1036
401 1036
2 1 17 0 0 8320 0 31 30 0 0 4
447 213
456 213
456 225
460 225
3 1 18 0 0 4224 0 32 31 0 0 2
387 213
411 213
2 0 19 0 0 4096 0 30 0 0 72 4
460 243
107 243
107 242
92 242
2 0 19 0 0 4096 0 7 0 0 72 2
455 1082
92 1082
3 2 20 0 0 4224 0 9 8 0 0 2
387 1054
401 1054
2 0 13 0 0 0 0 9 0 0 70 4
338 1063
238 1063
238 1062
223 1062
1 0 21 0 0 4096 0 9 0 0 71 2
338 1045
159 1045
3 2 22 0 0 8320 0 12 11 0 0 4
444 934
448 934
448 906
456 906
3 1 23 0 0 4224 0 14 11 0 0 3
441 854
441 888
456 888
2 0 21 0 0 4096 0 12 0 0 71 4
399 943
174 943
174 942
159 942
1 0 24 0 0 4096 0 13 0 0 62 2
341 889
249 889
2 0 19 0 0 0 0 14 0 0 72 2
395 863
92 863
1 3 25 0 0 8320 0 14 15 0 0 4
395 845
388 845
388 820
389 820
2 0 12 0 0 4096 0 15 0 0 61 2
344 829
315 829
1 0 24 0 0 4096 0 15 0 0 62 2
344 811
249 811
3 1 26 0 0 8320 0 17 16 0 0 3
389 729
389 742
457 742
2 0 27 0 0 4096 0 17 0 0 63 4
343 738
199 738
199 737
184 737
1 0 13 0 0 4096 0 17 0 0 70 2
343 720
223 720
2 0 12 0 0 4096 0 16 0 0 61 2
457 760
315 760
3 4 28 0 0 4224 0 18 19 0 0 4
489 602
397 602
397 652
385 652
1 3 29 0 0 8320 0 18 21 0 0 4
489 584
487 584
487 562
488 562
3 0 30 0 0 4096 0 19 0 0 69 2
340 661
287 661
2 0 24 0 0 0 0 19 0 0 62 4
340 652
264 652
264 653
249 653
1 0 21 0 0 0 0 19 0 0 71 4
340 643
174 643
174 642
159 642
2 0 12 0 0 0 0 20 0 0 61 2
338 614
315 614
1 0 13 0 0 0 0 20 0 0 70 2
338 596
223 596
2 0 27 0 0 4096 0 21 0 0 63 2
443 571
184 571
1 3 31 0 0 4224 0 21 22 0 0 3
443 553
443 545
435 545
2 0 12 0 0 0 0 22 0 0 61 2
389 554
315 554
2 0 13 0 0 0 0 23 0 0 70 2
340 525
223 525
1 0 19 0 0 0 0 23 0 0 72 2
340 507
92 507
2 0 30 0 0 4096 0 24 0 0 69 4
448 464
302 464
302 463
287 463
1 3 32 0 0 4224 0 24 25 0 0 4
448 446
399 446
399 424
386 424
2 0 24 0 0 0 0 25 0 0 62 4
340 433
264 433
264 432
249 432
1 0 21 0 0 0 0 25 0 0 71 2
340 415
159 415
2 0 27 0 0 4096 0 26 0 0 63 2
446 364
184 364
2 1 33 0 0 4224 0 27 26 0 0 3
441 320
441 346
446 346
1 3 34 0 0 4224 0 27 28 0 0 2
405 320
388 320
2 0 30 0 0 0 0 28 0 0 69 2
339 329
287 329
1 0 13 0 0 0 0 28 0 0 70 2
339 311
223 311
2 0 13 0 0 4096 0 29 0 0 70 4
523 262
305 262
305 263
223 263
3 1 35 0 0 8320 0 30 29 0 0 3
506 234
506 244
523 244
2 0 30 0 0 0 0 32 0 0 69 4
338 222
302 222
302 223
287 223
1 0 21 0 0 0 0 32 0 0 71 4
338 204
174 204
174 205
159 205
2 0 12 0 0 4224 0 33 0 0 0 2
315 171
315 1096
2 0 24 0 0 4224 0 34 0 0 0 2
249 174
249 1096
2 0 27 0 0 4224 0 35 0 0 0 2
184 172
184 1093
2 0 36 0 0 4224 0 36 0 0 0 2
119 172
119 1092
1 1 30 0 0 0 0 3 33 0 0 3
287 133
287 135
315 135
1 1 13 0 0 0 0 1 34 0 0 3
222 135
249 135
249 138
1 1 21 0 0 0 0 2 35 0 0 3
159 134
159 136
184 136
1 1 19 0 0 0 0 4 36 0 0 3
92 134
92 136
119 136
1 0 30 0 0 4224 0 3 0 0 0 2
287 133
287 1096
1 0 13 0 0 12416 0 1 0 0 0 4
222 135
222 263
223 263
223 1093
1 0 21 0 0 4224 0 2 0 0 0 2
159 134
159 1093
1 0 19 0 0 4224 0 4 0 0 0 2
92 134
92 1090
11
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
642 1051 678 1086
653 1059 666 1082
1 g
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
642 880 678 915
653 888 666 911
1 f
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
642 731 678 766
653 739 666 762
1 e
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
646 572 682 607
657 580 670 603
1 d
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
645 433 681 468
656 441 669 464
1 c
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
640 334 676 369
651 342 664 365
1 b
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
637 229 673 264
648 237 661 260
1 a
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
78 50 108 85
86 58 99 81
1 A
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
273 50 307 85
283 58 296 81
1 D
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
209 50 243 85
219 58 232 81
1 C
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
142 49 176 84
152 57 165 80
1 B
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
