CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
176 80 1364 707
110100498 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 255 60 0 1 11
0 24
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6369 0 0
2
43486.4 0
0
13 Logic Switch~
5 186 61 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9172 0 0
2
43486.4 0
0
13 Logic Switch~
5 127 60 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7100 0 0
2
43486.4 0
0
13 Logic Switch~
5 64 61 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3820 0 0
2
43486.4 0
0
7 Ground~
168 904 78 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7678 0 0
2
43486.5 0
0
8 2-In OR~
219 570 680 0 3 22
0 5 6 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
961 0 0
2
43486.5 0
0
8 2-In OR~
219 466 689 0 3 22
0 9 7 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
3178 0 0
2
43486.5 0
0
9 2-In AND~
219 368 710 0 3 22
0 8 3 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3409 0 0
2
43486.5 0
0
6 74136~
219 360 668 0 3 22
0 10 8 9
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3951 0 0
2
43486.5 0
0
8 2-In OR~
219 565 586 0 3 22
0 13 12 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
8885 0 0
2
43486.5 0
0
9 2-In AND~
219 464 621 0 3 22
0 14 10 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3780 0 0
2
43486.5 0
0
8 2-In OR~
219 359 612 0 3 22
0 15 3 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
9265 0 0
2
43486.5 0
0
8 2-In OR~
219 454 558 0 3 22
0 16 5 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
9442 0 0
2
43486.5 0
0
9 2-In AND~
219 368 549 0 3 22
0 15 3 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9424 0 0
2
43486.5 0
0
9 2-In AND~
219 447 497 0 3 22
0 18 3 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9968 0 0
2
43486.5 0
0
8 2-In OR~
219 356 488 0 3 22
0 19 8 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9281 0 0
2
43486.5 0
0
8 3-In OR~
219 568 385 0 4 22
0 23 22 21 20
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
8464 0 0
2
43486.5 0
0
5 7415~
219 365 432 0 4 22
0 10 15 24 21
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
7168 0 0
2
43486.5 0
0
9 2-In AND~
219 363 386 0 3 22
0 8 3 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3171 0 0
2
43486.4 0
0
9 2-In AND~
219 509 342 0 3 22
0 25 19 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4139 0 0
2
43486.4 0
0
8 2-In OR~
219 425 332 0 3 22
0 26 3 25
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
6435 0 0
2
43486.4 0
0
8 2-In OR~
219 352 324 0 3 22
0 5 8 26
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
5283 0 0
2
43486.4 0
0
8 2-In OR~
219 444 280 0 3 22
0 28 24 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6874 0 0
2
43486.4 0
0
8 2-In OR~
219 350 271 0 3 22
0 10 15 28
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
5305 0 0
2
43486.4 0
0
8 2-In OR~
219 499 229 0 3 22
0 30 19 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
34 0 0
2
43486.4 0
0
9 Inverter~
13 437 220 0 2 22
0 31 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
969 0 0
2
43486.4 0
0
6 74136~
219 373 220 0 3 22
0 8 24 31
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8402 0 0
2
43486.4 0
0
9 CC 7-Seg~
183 757 96 0 17 19
10 32 29 27 20 17 11 4 37 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
8 YELLOWCC
6 -41 62 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3751 0 0
2
43486.4 0
0
8 2-In OR~
219 588 183 0 3 22
0 33 8 32
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4292 0 0
2
43486.4 0
0
8 2-In OR~
219 503 174 0 3 22
0 34 5 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6118 0 0
2
43486.4 0
0
9 Inverter~
13 447 165 0 2 22
0 35 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
34 0 0
2
43486.4 0
0
6 74136~
219 372 165 0 3 22
0 10 24 35
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6357 0 0
2
43486.4 0
0
9 Inverter~
13 289 118 0 2 22
0 24 3
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
319 0 0
2
43486.4 0
0
9 Inverter~
13 220 118 0 2 22
0 8 15
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3976 0 0
2
43486.4 0
0
9 Inverter~
13 156 119 0 2 22
0 10 19
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7634 0 0
2
43486.4 0
0
9 Inverter~
13 90 116 0 2 22
0 5 36
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
523 0 0
2
43486.4 0
0
72
2 0 3 0 0 4096 0 21 0 0 7 2
412 341
292 341
2 0 3 0 0 0 0 19 0 0 7 2
339 395
292 395
2 0 3 0 0 4096 0 15 0 0 7 2
423 506
292 506
2 0 3 0 0 0 0 14 0 0 7 2
344 558
292 558
2 0 3 0 0 0 0 12 0 0 7 2
346 621
292 621
2 0 3 0 0 0 0 8 0 0 7 2
344 719
292 719
2 0 3 0 0 4224 0 33 0 0 0 2
292 136
292 742
3 7 4 0 0 8320 0 6 28 0 0 3
603 680
772 680
772 132
9 1 2 0 0 8320 0 28 5 0 0 4
757 54
757 29
904 29
904 72
1 0 5 0 0 12288 0 6 0 0 72 4
557 671
499 671
499 644
64 644
3 2 6 0 0 4224 0 7 6 0 0 2
499 689
557 689
3 2 7 0 0 4224 0 8 7 0 0 4
389 710
436 710
436 698
453 698
1 0 8 0 0 4096 0 8 0 0 68 2
344 701
186 701
3 1 9 0 0 4224 0 9 7 0 0 4
393 668
436 668
436 680
453 680
2 0 8 0 0 0 0 9 0 0 68 2
344 677
186 677
1 0 10 0 0 4096 0 9 0 0 70 2
344 659
127 659
3 6 11 0 0 8320 0 10 28 0 0 3
598 586
766 586
766 132
3 2 12 0 0 4224 0 11 10 0 0 4
485 621
520 621
520 595
552 595
3 1 13 0 0 4224 0 13 10 0 0 4
487 558
520 558
520 577
552 577
1 3 14 0 0 4224 0 11 12 0 0 2
440 612
392 612
2 0 10 0 0 4096 0 11 0 0 70 2
440 630
127 630
1 0 15 0 0 4096 0 12 0 0 67 2
346 603
223 603
1 3 16 0 0 4224 0 13 14 0 0 2
441 549
389 549
2 0 5 0 0 0 0 13 0 0 72 2
441 567
64 567
1 0 15 0 0 0 0 14 0 0 67 2
344 540
223 540
3 5 17 0 0 8320 0 15 28 0 0 3
468 497
760 497
760 132
1 3 18 0 0 4224 0 15 16 0 0 2
423 488
389 488
2 0 8 0 0 0 0 16 0 0 68 2
343 497
186 497
1 0 19 0 0 4096 0 16 0 0 69 2
343 479
159 479
4 4 20 0 0 8320 0 17 28 0 0 3
601 385
754 385
754 132
4 3 21 0 0 8320 0 18 17 0 0 3
386 432
386 394
555 394
3 2 22 0 0 8320 0 19 17 0 0 3
384 386
384 385
556 385
3 1 23 0 0 4224 0 20 17 0 0 3
530 342
530 376
555 376
3 0 24 0 0 4096 0 18 0 0 66 2
341 441
255 441
2 0 15 0 0 0 0 18 0 0 67 2
341 432
223 432
1 0 10 0 0 0 0 18 0 0 70 2
341 423
127 423
1 0 8 0 0 0 0 19 0 0 68 2
339 377
186 377
2 0 19 0 0 4096 0 20 0 0 69 2
485 351
159 351
3 1 25 0 0 8320 0 21 20 0 0 3
458 332
458 333
485 333
3 1 26 0 0 8320 0 22 21 0 0 3
385 324
385 323
412 323
2 0 8 0 0 0 0 22 0 0 68 2
339 333
186 333
1 0 5 0 0 0 0 22 0 0 72 2
339 315
64 315
3 3 27 0 0 4224 0 23 28 0 0 3
477 280
748 280
748 132
2 0 24 0 0 4096 0 23 0 0 66 2
431 289
255 289
1 3 28 0 0 4224 0 23 24 0 0 2
431 271
383 271
2 0 15 0 0 0 0 24 0 0 67 2
337 280
223 280
1 0 10 0 0 0 0 24 0 0 70 2
337 262
127 262
1 0 8 0 0 4096 0 27 0 0 68 2
357 211
186 211
3 2 29 0 0 4224 0 25 28 0 0 3
532 229
742 229
742 132
2 0 19 0 0 4096 0 25 0 0 69 2
486 238
159 238
2 1 30 0 0 4224 0 26 25 0 0 2
458 220
486 220
1 3 31 0 0 4224 0 26 27 0 0 2
422 220
406 220
2 0 24 0 0 0 0 27 0 0 66 2
357 229
255 229
3 1 32 0 0 4224 0 29 28 0 0 3
621 183
736 183
736 132
2 0 8 0 0 4096 0 29 0 0 68 2
575 192
186 192
3 1 33 0 0 4224 0 30 29 0 0 2
536 174
575 174
2 0 5 0 0 128 0 30 0 0 72 2
490 183
64 183
2 1 34 0 0 4224 0 31 30 0 0 2
468 165
490 165
3 1 35 0 0 4224 0 32 31 0 0 2
405 165
432 165
2 0 24 0 0 0 0 32 0 0 66 2
356 174
255 174
1 0 10 0 0 0 0 32 0 0 70 2
356 156
127 156
1 0 24 0 0 0 0 33 0 0 66 3
292 100
292 77
255 77
1 0 8 0 0 0 0 34 0 0 68 3
223 100
223 77
186 77
1 0 10 0 0 0 0 35 0 0 70 3
159 101
159 77
127 77
1 0 5 0 0 0 0 36 0 0 72 3
93 98
93 78
64 78
1 0 24 0 0 4224 0 1 0 0 0 2
255 72
255 721
2 0 15 0 0 4224 0 34 0 0 0 2
223 136
223 721
1 0 8 0 0 4224 0 2 0 0 0 2
186 73
186 720
2 0 19 0 0 4224 0 35 0 0 0 2
159 137
159 720
1 0 10 0 0 4224 0 3 0 0 0 2
127 72
127 721
2 0 36 0 0 4224 0 36 0 0 0 2
93 134
93 720
1 0 5 0 0 4224 0 4 0 0 0 2
64 73
64 721
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
