CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 225 59 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 162 59 0 1 11
0 18
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89878e-315 5.26354e-315
0
13 Logic Switch~
5 107 60 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89878e-315 5.30499e-315
0
13 Logic Switch~
5 52 57 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89878e-315 5.32571e-315
0
10 2-In XNOR~
219 268 130 0 3 22
0 5 4 3
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
8157 0 0
2
43490.4 0
0
8 2-In OR~
219 383 235 0 3 22
0 7 8 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
5572 0 0
2
5.89878e-315 5.34643e-315
0
9 Inverter~
13 316 204 0 2 22
0 9 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
8901 0 0
2
5.89878e-315 5.3568e-315
0
9 2-In XOR~
219 270 204 0 3 22
0 18 4 9
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7361 0 0
2
5.89878e-315 5.36716e-315
0
8 3-In OR~
219 341 167 0 4 22
0 3 13 18 10
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U11B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 11 0
1 U
4747 0 0
2
5.89878e-315 5.37752e-315
0
8 3-In OR~
219 399 632 0 4 22
0 13 12 15 14
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U11A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 11 0
1 U
972 0 0
2
5.89878e-315 5.38788e-315
0
9 2-In AND~
219 283 605 0 3 22
0 17 16 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3472 0 0
2
5.89878e-315 5.39306e-315
0
9 Inverter~
13 238 92 0 2 22
0 4 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9998 0 0
2
5.89878e-315 5.39824e-315
0
9 2-In AND~
219 343 357 0 3 22
0 24 8 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3536 0 0
2
5.89878e-315 5.40342e-315
0
7 Ground~
168 805 156 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.89878e-315 5.4086e-315
0
8 3-In OR~
219 344 771 0 4 22
0 30 31 13 26
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 7 0
1 U
3835 0 0
2
5.89878e-315 5.41378e-315
0
9 2-In XOR~
219 278 771 0 3 22
0 5 18 31
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3670 0 0
2
5.89878e-315 5.41896e-315
0
9 2-In AND~
219 284 726 0 3 22
0 16 18 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
5616 0 0
2
5.89878e-315 5.42414e-315
0
9 2-In AND~
219 344 690 0 3 22
0 19 5 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9323 0 0
2
5.89878e-315 5.42933e-315
0
8 2-In OR~
219 274 654 0 3 22
0 17 16 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
317 0 0
2
5.89878e-315 5.43192e-315
0
9 2-In AND~
219 349 518 0 3 22
0 20 16 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3108 0 0
2
5.89878e-315 5.43451e-315
0
8 2-In OR~
219 273 485 0 3 22
0 8 18 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4299 0 0
2
5.89878e-315 5.4371e-315
0
8 3-In OR~
219 400 409 0 4 22
0 21 23 22 28
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
9672 0 0
2
5.89878e-315 5.43969e-315
0
5 7415~
219 284 438 0 4 22
0 5 17 4 22
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
7876 0 0
2
5.89878e-315 5.44228e-315
0
9 2-In AND~
219 283 393 0 3 22
0 18 16 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
6369 0 0
2
5.89878e-315 5.44487e-315
0
8 3-In OR~
219 276 321 0 4 22
0 13 18 16 24
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 3 0
1 U
9172 0 0
2
5.89878e-315 5.44746e-315
0
8 3-In OR~
219 275 278 0 4 22
0 5 17 4 29
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 3 0
1 U
7100 0 0
2
5.89878e-315 5.45005e-315
0
9 Inverter~
13 174 94 0 2 22
0 18 17
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3820 0 0
2
5.89878e-315 5.45264e-315
0
9 Inverter~
13 121 94 0 2 22
0 5 8
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7678 0 0
2
5.89878e-315 5.45523e-315
0
9 Inverter~
13 67 96 0 2 22
0 13 25
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
961 0 0
2
5.89878e-315 5.45782e-315
0
9 CC 7-Seg~
183 705 95 0 17 19
10 10 6 29 28 27 14 26 32 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3178 0 0
2
5.89878e-315 5.46041e-315
0
79
3 0 3 0 0 0 0 5 0 0 4 2
307 130
307 130
2 0 4 0 0 4096 0 8 0 0 56 2
254 213
225 213
1 0 5 0 0 4096 0 5 0 0 59 2
252 121
107 121
0 1 3 0 0 8320 0 0 9 0 0 4
302 130
313 130
313 158
328 158
3 2 6 0 0 4224 0 6 30 0 0 3
416 235
690 235
690 131
2 1 7 0 0 8320 0 7 6 0 0 4
337 204
357 204
357 226
370 226
2 0 8 0 0 4096 0 6 0 0 62 2
370 244
124 244
1 3 9 0 0 4224 0 7 8 0 0 2
301 204
303 204
4 0 10 0 0 0 0 9 0 0 69 2
374 167
374 167
0 0 11 0 0 8320 0 0 0 0 0 3
297 129
297 130
302 130
3 2 12 0 0 12416 0 11 10 0 0 4
304 605
320 605
320 632
387 632
0 1 13 0 0 4096 0 0 10 61 0 4
52 578
371 578
371 623
386 623
4 0 14 0 0 8192 0 10 0 0 65 3
432 632
432 631
435 631
3 0 15 0 0 8192 0 10 0 0 29 3
386 641
386 640
382 640
2 0 16 0 0 4096 0 11 0 0 22 2
259 614
241 614
1 0 17 0 0 4096 0 11 0 0 58 2
259 596
177 596
1 0 16 0 0 4096 0 17 0 0 22 2
260 717
241 717
2 0 16 0 0 4096 0 19 0 0 22 2
261 663
241 663
2 0 16 0 0 4096 0 20 0 0 22 2
325 527
241 527
2 0 16 0 0 0 0 24 0 0 22 2
259 402
241 402
3 0 16 0 0 0 0 25 0 0 22 2
263 330
241 330
2 0 16 0 0 4224 0 12 0 0 0 2
241 110
241 900
2 0 13 0 0 0 0 9 0 0 61 2
329 167
52 167
1 0 5 0 0 0 0 28 0 0 59 2
124 76
107 76
1 0 18 0 0 4096 0 27 0 0 57 2
177 76
162 76
1 0 4 0 0 0 0 12 0 0 56 3
241 74
241 75
225 75
0 1 13 0 0 0 0 0 29 61 0 3
52 76
52 78
70 78
3 1 19 0 0 8320 0 19 18 0 0 3
307 654
320 654
320 681
3 3 15 0 0 12416 0 10 18 0 0 5
386 641
386 640
369 640
369 690
365 690
2 0 18 0 0 4096 0 21 0 0 57 2
260 494
162 494
3 1 20 0 0 8320 0 21 20 0 0 4
306 485
319 485
319 509
325 509
3 1 21 0 0 8320 0 13 22 0 0 4
364 357
372 357
372 400
387 400
3 4 22 0 0 12416 0 22 23 0 0 4
387 418
349 418
349 438
305 438
3 2 23 0 0 4224 0 24 22 0 0 4
304 393
348 393
348 409
388 409
3 0 4 0 0 4096 0 23 0 0 56 2
260 447
225 447
2 0 17 0 0 4096 0 23 0 0 58 2
260 438
177 438
1 0 5 0 0 4096 0 23 0 0 59 2
260 429
107 429
1 0 18 0 0 0 0 24 0 0 57 2
259 384
162 384
3 0 13 0 0 0 0 15 0 0 61 4
331 780
327 780
327 793
52 793
2 0 18 0 0 4096 0 16 0 0 57 2
262 780
162 780
1 0 5 0 0 4096 0 16 0 0 59 2
262 762
107 762
2 0 18 0 0 0 0 17 0 0 57 2
260 735
162 735
2 0 5 0 0 4096 0 18 0 0 59 2
320 699
107 699
1 0 17 0 0 4096 0 19 0 0 58 2
261 645
177 645
1 0 8 0 0 0 0 21 0 0 62 2
260 476
124 476
2 0 8 0 0 0 0 13 0 0 62 2
319 366
124 366
4 1 24 0 0 8320 0 25 13 0 0 4
309 321
313 321
313 348
319 348
2 0 18 0 0 4096 0 25 0 0 57 2
264 321
162 321
1 0 13 0 0 0 0 25 0 0 61 2
263 312
52 312
1 0 18 0 0 0 0 8 0 0 57 2
254 195
162 195
1 0 5 0 0 0 0 26 0 0 59 2
262 269
107 269
2 0 17 0 0 4096 0 26 0 0 58 2
263 278
177 278
3 0 4 0 0 4096 0 26 0 0 56 2
262 287
225 287
3 0 18 0 0 4096 0 9 0 0 57 2
328 176
162 176
2 0 4 0 0 0 0 5 0 0 56 2
252 139
225 139
1 0 4 0 0 4224 0 1 0 0 0 2
225 71
225 891
1 0 18 0 0 4224 0 2 0 0 0 2
162 71
162 880
2 0 17 0 0 4224 0 27 0 0 0 2
177 112
177 891
1 0 5 0 0 4224 0 3 0 0 0 2
107 72
107 897
2 0 25 0 0 4224 0 29 0 0 0 2
70 114
70 900
1 0 13 0 0 4224 0 4 0 0 0 2
52 69
52 900
2 0 8 0 0 4224 0 28 0 0 0 2
124 112
124 899
9 1 2 0 0 12416 0 30 14 0 0 4
705 53
705 23
805 23
805 150
7 4 26 0 0 4224 0 30 15 0 0 3
720 131
720 771
377 771
4 6 14 0 0 12416 0 10 30 0 0 4
432 632
432 631
714 631
714 131
3 5 27 0 0 8320 0 20 30 0 0 3
370 518
708 518
708 131
4 4 28 0 0 8320 0 22 30 0 0 3
433 409
702 409
702 131
4 3 29 0 0 4224 0 26 30 0 0 3
308 278
696 278
696 131
0 1 10 0 0 4224 0 0 30 0 0 3
371 167
684 167
684 131
3 1 30 0 0 8320 0 17 15 0 0 4
305 726
326 726
326 762
331 762
3 2 31 0 0 4224 0 16 15 0 0 2
311 771
332 771
3 3 4 0 0 0 0 23 23 0 0 2
260 447
260 447
2 2 17 0 0 0 0 23 23 0 0 2
260 438
260 438
1 1 5 0 0 0 0 23 23 0 0 2
260 429
260 429
2 2 16 0 0 0 0 24 24 0 0 2
259 402
259 402
1 1 18 0 0 0 0 24 24 0 0 2
259 384
259 384
3 3 4 0 0 0 0 26 26 0 0 2
262 287
262 287
2 2 17 0 0 0 0 26 26 0 0 2
263 278
263 278
1 1 5 0 0 0 0 26 26 0 0 2
262 269
262 269
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
